----------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

entity mario_easy is
port (
	clk		: in std_logic;     -- 25MHz
	p1       : in std_logic;
	rss      : in std_logic;
	note_clk : out std_logic;
	d_d      : out std_logic_vector(9 downto 0);
	d_dp     : out std_logic_vector(9 downto 0);
	d_dm     : out std_logic_vector(9 downto 0);	
	reset    : out std_logic;
	rr       : in std_logic;
   -------------------------------------------------------dot port
	dot_d : out std_logic_vector ( 9 downto 0);
	dot_scan : out std_logic_vector ( 13 downto 0);
	--------------------------------------------------------piezo port
	piezo	   : out std_logic;
	piezo2   : out std_logic;
	led : out std_logic
);
end mario_easy;

architecture a of mario_easy is
-------------------------------------------------------------------------------component
component dot_dis
port (
	clk : in std_logic;
	dot_data_00 : in std_logic_vector (9 downto 0);
	dot_data_01 : in std_logic_vector (9 downto 0);
	dot_data_02 : in std_logic_vector (9 downto 0);
	dot_data_03 : in std_logic_vector (9 downto 0);
	dot_data_04 : in std_logic_vector (9 downto 0);
	dot_data_05 : in std_logic_vector (9 downto 0);
	dot_data_06 : in std_logic_vector (9 downto 0);
	dot_data_07 : in std_logic_vector (9 downto 0);
	dot_data_08 : in std_logic_vector (9 downto 0);
	dot_data_09 : in std_logic_vector (9 downto 0);
	dot_data_10 : in std_logic_vector (9 downto 0);
	dot_data_11 : in std_logic_vector (9 downto 0);
	dot_data_12 : in std_logic_vector (9 downto 0);
	dot_data_13 : in std_logic_vector (9 downto 0);

	dot_d : out std_logic_vector (9 downto 0);
	dot_scan : out std_logic_vector ( 13 downto 0)
);
end component;
------------------------------------------------------------------------com signal
signal ryt  : integer range 0 to 920312;
signal note : integer range 0 to 1500 := 1450;
signal n_clk   : std_logic := '0';
signal rst : std_logic := '0';

---------------------------------------------------------------------dot signal
signal dot_data_00 : std_logic_vector (9 downto 0);
signal dot_data_01 : std_logic_vector (9 downto 0);
signal dot_data_02 : std_logic_vector (9 downto 0);
signal dot_data_03 : std_logic_vector (9 downto 0);
signal dot_data_04 : std_logic_vector (9 downto 0);
signal dot_data_05 : std_logic_vector (9 downto 0);
signal dot_data_06 : std_logic_vector (9 downto 0);
signal dot_data_07 : std_logic_vector (9 downto 0);
signal dot_data_08 : std_logic_vector (9 downto 0);
signal dot_data_09 : std_logic_vector (9 downto 0);
signal dot_data_10 : std_logic_vector (9 downto 0);
signal dot_data_11 : std_logic_vector (9 downto 0);
signal dot_data_12 : std_logic_vector (9 downto 0);
signal dot_data_13 : std_logic_vector (9 downto 0);

constant zr : std_logic_vector(9 downto 0) := "0000000000";

type data_a is array(1500 downto 0) of std_logic_vector(9 downto 0);
signal data_b : data_a;

--------------------------------------------------------------------piezo signal
constant r  : integer range 0 to 1000000 := 0;

constant a_1 	: integer range 0 to 1000000 := 454544;
constant bm_1 	: integer range 0 to 1000000 := 429034;
constant b_1 	: integer range 0 to 1000000 := 404954;
constant c_1 	: integer range 0 to 1000000 := 382226;
constant dm_1 	: integer range 0 to 1000000 := 360773;
constant d_1 	: integer range 0 to 1000000 := 340524;
constant em_1 	: integer range 0 to 1000000 := 321414;
constant e_1 	: integer range 0 to 1000000 := 303373;
constant f_1 	: integer range 0 to 1000000 := 286346;
constant gm_1 	: integer range 0 to 1000000 := 270274;
constant g_1 	: integer range 0 to 1000000 := 255105;
constant am_1 	: integer range 0 to 1000000 := 240787;

constant a_2 	: integer range 0 to 1000000 := 227273;
constant bm_2 	: integer range 0 to 1000000 := 214517;
constant b_2 	: integer range 0 to 1000000 := 202477;
constant c_2 	: integer range 0 to 1000000 := 191113;
constant dm_2 	: integer range 0 to 1000000 := 180387;
constant d_2 	: integer range 0 to 1000000 := 170262;
constant em_2 	: integer range 0 to 1000000 := 160706;
constant e_2 	: integer range 0 to 1000000 := 151686;
constant f_2 	: integer range 0 to 1000000 := 143173;
constant gm_2 	: integer range 0 to 1000000 := 135137;
constant g_2 	: integer range 0 to 1000000 := 127553;
constant am_2 	: integer range 0 to 1000000 := 120394;

constant a_3 	: integer range 0 to 1000000 := 113635;
constant bm_3 	: integer range 0 to 1000000 := 107257;
constant b_3 	: integer range 0 to 1000000 := 101237;
constant c_3 	: integer range 0 to 1000000 := 95555;
constant dm_3 	: integer range 0 to 1000000 := 90192;
constant d_3 	: integer range 0 to 1000000 := 85130;
constant em_3 	: integer range 0 to 1000000 := 80352;
constant e_3 	: integer range 0 to 1000000 := 75842;
constant f_3 	: integer range 0 to 1000000 := 71585;
constant gm_3 	: integer range 0 to 1000000 := 67568;
constant g_3 	: integer range 0 to 1000000 := 63775;
constant am_3 	: integer range 0 to 1000000 := 60196;

constant a_4 	: integer range 0 to 1000000 := 56817;
constant bm_4 	: integer range 0 to 1000000 := 53628;
constant b_4 	: integer range 0 to 1000000 := 50618;
constant c_4 	: integer range 0 to 1000000 := 47777;
constant dm_4 	: integer range 0 to 1000000 := 45096;
constant d_4 	: integer range 0 to 1000000 := 42565;
constant em_4 	: integer range 0 to 1000000 := 40176;
constant e_4 	: integer range 0 to 1000000 := 37921;
constant f_4 	: integer range 0 to 1000000 := 35792;
constant gm_4 	: integer range 0 to 1000000 := 33783;
constant g_4 	: integer range 0 to 1000000 := 31887;
constant am_4 	: integer range 0 to 1000000 := 30097;

constant a_5 	: integer range 0 to 1000000 := 28408;
constant bm_5 	: integer range 0 to 1000000 := 26814;
constant b_5 	: integer range 0 to 1000000 := 25309;
constant c_5 	: integer range 0 to 1000000 := 23888;
constant dm_5 	: integer range 0 to 1000000 := 22547;
constant d_5 	: integer range 0 to 1000000 := 21282;
constant em_5 	: integer range 0 to 1000000 := 20087;
constant e_5 	: integer range 0 to 1000000 := 18960;
constant f_5 	: integer range 0 to 1000000 := 17896;
constant gm_5 	: integer range 0 to 1000000 := 16891;
constant g_5 	: integer range 0 to 1000000 := 15943;
constant am_5 	: integer range 0 to 1000000 := 15048;

constant a_6 	: integer range 0 to 1000000 := 14204;
constant bm_6 	: integer range 0 to 1000000 := 13406;
constant b_6 	: integer range 0 to 1000000 := 12654;
constant c_6 	: integer range 0 to 1000000 := 11945;
constant dm_6 	: integer range 0 to 1000000 := 11273;
constant d_6 	: integer range 0 to 1000000 := 10640;
constant em_6 	: integer range 0 to 1000000 := 10043;
constant e_6 	: integer range 0 to 1000000 := 9479;
constant f_6 	: integer range 0 to 1000000 := 8947;
constant gm_6 	: integer range 0 to 1000000 := 8445;
constant g_6 	: integer range 0 to 1000000 := 7971;
constant am_6 	: integer range 0 to 1000000 := 7524;


signal cnt 	: integer range 0 to 1000000;
signal cnt2 : integer range 0 to 1000000;
signal seq  : integer range 0 to 100000;


signal st   : std_logic := '0';

signal p_clk	: std_logic;
signal p_clk2  : std_logic;

type scale_a is array (1500 downto 0) of integer range 0 to 1000000;
signal scale : scale_a;
signal scale2: scale_a;
------------------------------------------------------------------------com

begin

process(p1,rss,rst)
begin
  if p1 = '1' then
     st <= '1';
  elsif rst = '1' or rss = '1' then
     st <= '0';
	  seq <= 0;
  end if;
end process;

process(clk,rst,rss)
begin
  if rst = '1' or rss = '1' then
     ryt <= 0;
	  n_clk <= '0';
  elsif clk'event and clk = '1' and st = '1' then
     if ryt = 920312 then
	     ryt <= 0;
        n_clk <= not n_clk;
     else
        ryt <= ryt + 1;
        n_clk <= n_clk;		  
     end if;
  end if;
end process;

note_clk <= n_clk;

process(n_clk,rss,rst,clk)
begin
  if rss = '1' or rst = '1' then
     note <= 1450;
  elsif n_clk'event and n_clk = '1' then
     if note = 1440 then
	     note <= 1450;
		  rst <= '1';
	  elsif note = 1500 then
	     note <= 0;
	  else
		  note <= note + 1;
     end if;
  end if;
  if rss = '1' or rr = '1' then
     rst <= '0';
  end if;  
end process;

reset <= rst;

---------------------------------------------------------------------dot
data_b(0) <= "0000000001";
data_b(1) <= "0000000000";
data_b(2) <= "0000000001";
data_b(3) <= "0000000000";
data_b(4) <= "0000000000";
data_b(5) <= "0000000000";
data_b(6) <= "0000000001";
data_b(7) <= "0000000000";
data_b(8) <= "0000000000";
data_b(9) <= "0000000000";
data_b(10) <= "0000000010";
data_b(11) <= "0000000000";
data_b(12) <= "0000000001";
data_b(13) <= "0000000000";
data_b(14) <= "0000000000";
data_b(15) <= "0000000000";
--------------------------------1
data_b(16) <= "0000000001";
data_b(17) <= "0000000000";
data_b(18) <= "0000000000";
data_b(19) <= "0000000000";
data_b(20) <= "0000000000";
data_b(21) <= "0000000000";
data_b(22) <= "0000000000";
data_b(23) <= "0000000000";
data_b(24) <= "0010000000";
data_b(25) <= "0000000000";
data_b(26) <= "0000000000";
data_b(27) <= "0000000000";
data_b(28) <= "0000000000";
data_b(29) <= "0000000000";
data_b(30) <= "0000000000";
data_b(31) <= "0000000000";
-----------------------------------2
data_b(32) <= "0000000010";
data_b(33) <= "0000000000";
data_b(34) <= "0000000000";
data_b(35) <= "0000000000";
data_b(36) <= "0000000000";
data_b(37) <= "0000000000";
data_b(38) <= "0000000100";
data_b(39) <= "0000000000";
data_b(40) <= "0000000000";
data_b(41) <= "0000000000";
data_b(42) <= "0000000000";
data_b(43) <= "0000000000";
data_b(44) <= "0010000000";
data_b(45) <= "0000000000";
data_b(46) <= "0000000000";
data_b(47) <= "0000000000";
----------------------------------3
data_b(48) <= "0000000000";
data_b(49) <= "0000000000";
data_b(50) <= "0000000100";
data_b(51) <= "0000000000";
data_b(52) <= "0000000000";
data_b(53) <= "0000000000";
data_b(54) <= "0000000010";
data_b(55) <= "0000000000";
data_b(56) <= "0000000000";
data_b(57) <= "0000000000";
data_b(58) <= "0000000010";
data_b(59) <= "0000000000";
data_b(60) <= "0000000100";
data_b(61) <= "0000000000";
data_b(62) <= "0000000000";
data_b(63) <= "0000000000";
-----------------------------------4
data_b(64) <= "0010000000";
data_b(65) <= "0000000000";
data_b(66) <= "0000000000";
data_b(67) <= "0000000100";
data_b(68) <= "0000000000";
data_b(69) <= "0000000000";
data_b(70) <= "0000000010";
data_b(71) <= "0000000000";
data_b(72) <= "0000000001";
data_b(73) <= "0000000000";
data_b(74) <= "0000000000";
data_b(75) <= "0000000000";
data_b(76) <= "0000000010";
data_b(77) <= "0000000000";
data_b(78) <= "0000000001";
data_b(79) <= "0000000000";
-----------------------------------5
data_b(80) <= "0000000000";
data_b(81) <= "0000000000";
data_b(82) <= "0000000001";
data_b(83) <= "0000000000";
data_b(84) <= "0000000000";
data_b(85) <= "0000000000";
data_b(86) <= "0000000100";
data_b(87) <= "0000000000";
data_b(88) <= "0000000010";
data_b(89) <= "0000000000";
data_b(90) <= "0010000000";
data_b(91) <= "0000000000";
data_b(92) <= "0000000000";
data_b(93) <= "0000000000";
data_b(94) <= "0000000000";
data_b(95) <= "0000000000";
------------------------------------6
data_b(96) <= "0000000001";
data_b(97) <= "0000000000";
data_b(98) <= "0000000000";
data_b(99) <= "0000000000";
data_b(100) <= "0000000000";
data_b(101) <= "0000000000";
data_b(102) <= "0000000010";
data_b(103) <= "0000000000";
data_b(104) <= "0000000000";
data_b(105) <= "0000000000";
data_b(106) <= "0000000000";
data_b(107) <= "0000000000";
data_b(108) <= "0000000100";
data_b(109) <= "0000000000";
data_b(110) <= "0000000000";
data_b(111) <= "0000000000";
----------------------------------7
data_b(112) <= "0000000000";
data_b(113) <= "0000000000";
data_b(114) <= "0100000000";
data_b(115) <= "0000000000";
data_b(116) <= "0000000000";
data_b(117) <= "0000000000";
data_b(118) <= "0010000000";
data_b(119) <= "0000000000";
data_b(120) <= "0000000000";
data_b(121) <= "0000000000";
data_b(122) <= "0010000000";
data_b(123) <= "0000000000";
data_b(124) <= "0100000000";
data_b(125) <= "0000000000";
data_b(126) <= "0000000000";
data_b(127) <= "0000000000";
-----------------------------------8
data_b(128) <= "0010000000";
data_b(129) <= "0000000000";
data_b(130) <= "0000000000";
data_b(131) <= "0000000100";
data_b(132) <= "0000000000";
data_b(133) <= "0000000000";
data_b(134) <= "0000000010";
data_b(135) <= "0000000000";
data_b(136) <= "0000000001";
data_b(137) <= "0000000000";
data_b(138) <= "0000000000";
data_b(139) <= "0000000000";
data_b(140) <= "0000000010";
data_b(141) <= "0000000000";
data_b(142) <= "0000000001";
data_b(143) <= "0000000000";
-----------------------------------9
data_b(144) <= "0000000000";
data_b(145) <= "0000000000";
data_b(146) <= "0000000001";
data_b(147) <= "0000000000";
data_b(148) <= "0000000000";
data_b(149) <= "0000000000";
data_b(150) <= "0000000100";
data_b(151) <= "0000000000";
data_b(152) <= "0000000010";
data_b(153) <= "0000000000";
data_b(154) <= "0010000000";
data_b(155) <= "0000000000";
data_b(156) <= "0000000000";
data_b(157) <= "0000000000";
data_b(158) <= "0000000000";
data_b(159) <= "0000000000";
------------------------------------10
data_b(160) <= "0000000000";
data_b(161) <= "0000000000";
data_b(162) <= "0000000000";
data_b(163) <= "0000000000";
data_b(164) <= "0000000001";
data_b(165) <= "0000000000";
data_b(166) <= "0000000010";
data_b(167) <= "0000000000";
data_b(168) <= "0000000010";
data_b(169) <= "0000000000";
data_b(170) <= "0010000000";
data_b(171) <= "0000000000";
data_b(172) <= "0000000000";
data_b(173) <= "0000000000";
data_b(174) <= "0000000010";
data_b(175) <= "0000000000";
--------------------------------11
data_b(176) <= "0000000000";
data_b(177) <= "0000000000";
data_b(178) <= "0010000000";
data_b(179) <= "0000000000";
data_b(180) <= "0000000100";
data_b(181) <= "0000000000";
data_b(182) <= "0000000010";
data_b(183) <= "0000000000";
data_b(184) <= "0000000000";
data_b(185) <= "0000000000";
data_b(186) <= "0000000100";
data_b(187) <= "0000000000";
data_b(188) <= "0000000010";
data_b(189) <= "0000000000";
data_b(190) <= "0000000001";
data_b(191) <= "0000000000";
----------------------------------12
data_b(192) <= "0000000000";
data_b(193) <= "0000000000";
data_b(194) <= "0000000000";
data_b(195) <= "0000000000";
data_b(196) <= "0000000001";
data_b(197) <= "0000000000";
data_b(198) <= "0000000010";
data_b(199) <= "0000000000";
data_b(200) <= "0000000010";
data_b(201) <= "0000000000";
data_b(202) <= "0000000100";
data_b(203) <= "0000000000";
data_b(204) <= "0000000000";
data_b(205) <= "0000000000";
data_b(206) <= "0000000010";
data_b(207) <= "0000000000";
--------------------------------13
data_b(208) <= "0000000000";
data_b(209) <= "0000000000";
data_b(210) <= "1000000000";
data_b(211) <= "0000000000";
data_b(212) <= "0000000000";
data_b(213) <= "0000000000";
data_b(214) <= "1000000000";
data_b(215) <= "0000000000";
data_b(216) <= "1000000000";
data_b(217) <= "0000000000";
data_b(218) <= "0000000000";
data_b(219) <= "0000000000";
data_b(220) <= "0000000100";
data_b(221) <= "0000000000";
data_b(222) <= "0000000000";
data_b(223) <= "0000000000";
-------------------------------14
data_b(224) <= "0000000000";
data_b(225) <= "0000000000";
data_b(226) <= "0000000000";
data_b(227) <= "0000000000";
data_b(228) <= "0000000001";
data_b(229) <= "0000000000";
data_b(230) <= "0000000010";
data_b(231) <= "0000000000";
data_b(232) <= "0000000010";
data_b(233) <= "0000000000";
data_b(234) <= "0000000100";
data_b(235) <= "0000000000";
data_b(236) <= "0000000000";
data_b(237) <= "0000000000";
data_b(238) <= "0000000010";
data_b(239) <= "0000000000";
-------------------------------15
data_b(240) <= "0000000000";
data_b(241) <= "0000000000";
data_b(242) <= "0010000000";
data_b(243) <= "0000000000";
data_b(244) <= "0000000100";
data_b(245) <= "0000000000";
data_b(246) <= "0000000010";
data_b(247) <= "0000000000";
data_b(248) <= "0000000000";
data_b(249) <= "0000000000";
data_b(250) <= "0000000100";
data_b(251) <= "0000000000";
data_b(252) <= "0000000010";
data_b(253) <= "0000000000";
data_b(254) <= "0000000001";
data_b(255) <= "0000000000";
-----------------------------16
data_b(256) <= "0000000000";
data_b(257) <= "0000000000";
data_b(258) <= "0000000000";
data_b(259) <= "0000000000";
data_b(260) <= "0100000000";
data_b(261) <= "0000000000";
data_b(262) <= "0000000000";
data_b(263) <= "0000000000";
data_b(264) <= "0000000000";
data_b(265) <= "0000000000";
data_b(266) <= "0010000000";
data_b(267) <= "0000000000";
data_b(268) <= "0000000000";
data_b(269) <= "0000000000";
data_b(270) <= "0000000000";
data_b(271) <= "0000000000";
-------------------------------17
data_b(272) <= "0000000100";
data_b(273) <= "0000000000";
data_b(274) <= "0000000000";
data_b(275) <= "0000000000";
data_b(276) <= "0000000000";
data_b(277) <= "0000000000";
data_b(278) <= "0010000000";
data_b(279) <= "0000000000";
data_b(280) <= "0010000000";
data_b(281) <= "0000000000";
data_b(282) <= "0000000000";
data_b(283) <= "0000000000";
data_b(284) <= "1000000000";
data_b(285) <= "0000000000";
data_b(286) <= "0000000000";
data_b(287) <= "0000000000";
--------------------------------18
data_b(288) <= "0000000000";
data_b(289) <= "0000000000";
data_b(290) <= "0000000000";
data_b(291) <= "0000000000";
data_b(292) <= "0000000001";
data_b(293) <= "0000000000";
data_b(294) <= "0000000010";
data_b(295) <= "0000000000";
data_b(296) <= "0000000010";
data_b(297) <= "0000000000";
data_b(298) <= "0010000000";
data_b(299) <= "0000000000";
data_b(300) <= "0000000000";
data_b(301) <= "0000000000";
data_b(302) <= "0000000010";
data_b(303) <= "0000000000";
-------------------------------19
data_b(304) <= "0000000000";
data_b(305) <= "0000000000";
data_b(306) <= "0010000000";
data_b(307) <= "0000000000";
data_b(308) <= "0000000100";
data_b(309) <= "0000000000";
data_b(310) <= "0000000010";
data_b(311) <= "0000000000";
data_b(312) <= "0000000000";
data_b(313) <= "0000000000";
data_b(314) <= "0000000100";
data_b(315) <= "0000000000";
data_b(316) <= "0000000010";
data_b(317) <= "0000000000";
data_b(318) <= "0000000001";
data_b(319) <= "0000000000";
----------------------------------20
data_b(320) <= "0000000000";
data_b(321) <= "0000000000";
data_b(322) <= "0000000000";
data_b(323) <= "0000000000";
data_b(324) <= "0000000001";
data_b(325) <= "0000000000";
data_b(326) <= "0000000010";
data_b(327) <= "0000000000";
data_b(328) <= "0000000010";
data_b(329) <= "0000000000";
data_b(330) <= "0000000100";
data_b(331) <= "0000000000";
data_b(332) <= "0000000000";
data_b(333) <= "0000000000";
data_b(334) <= "0000000010";
data_b(335) <= "0000000000";
--------------------------------21
data_b(336) <= "0000000000";
data_b(337) <= "0000000000";
data_b(338) <= "1000000000";
data_b(339) <= "0000000000";
data_b(340) <= "0000000000";
data_b(341) <= "0000000000";
data_b(342) <= "1000000000";
data_b(343) <= "0000000000";
data_b(344) <= "1000000000";
data_b(345) <= "0000000000";
data_b(346) <= "0000000000";
data_b(347) <= "0000000000";
data_b(348) <= "0000000100";
data_b(349) <= "0000000000";
data_b(350) <= "0000000000";
data_b(351) <= "0000000000";
---------------------------------22
data_b(352) <= "0000000000";
data_b(353) <= "0000000000";
data_b(354) <= "0000000000";
data_b(355) <= "0000000000";
data_b(356) <= "0000000001";
data_b(357) <= "0000000000";
data_b(358) <= "0000000010";
data_b(359) <= "0000000000";
data_b(360) <= "0000000010";
data_b(361) <= "0000000000";
data_b(362) <= "0000000100";
data_b(363) <= "0000000000";
data_b(364) <= "0000000000";
data_b(365) <= "0000000000";
data_b(366) <= "0000000010";
data_b(367) <= "0000000000";
------------------------------23
data_b(368) <= "0000000000";
data_b(369) <= "0000000000";
data_b(370) <= "0010000000";
data_b(371) <= "0000000000";
data_b(372) <= "0000000100";
data_b(373) <= "0000000000";
data_b(374) <= "0000000010";
data_b(375) <= "0000000000";
data_b(376) <= "0000000000";
data_b(377) <= "0000000000";
data_b(378) <= "0000000100";
data_b(379) <= "0000000000";
data_b(380) <= "0000000010";
data_b(381) <= "0000000000";
data_b(382) <= "0000000001";
data_b(383) <= "0000000000";
----------------------------24
data_b(384) <= "0000000000";
data_b(385) <= "0000000000";
data_b(386) <= "0000000000";
data_b(387) <= "0000000000";
data_b(388) <= "0100000000";
data_b(389) <= "0000000000";
data_b(390) <= "0000000000";
data_b(391) <= "0000000000";
data_b(392) <= "0000000000";
data_b(393) <= "0000000000";
data_b(394) <= "0010000000";
data_b(395) <= "0000000000";
data_b(396) <= "0000000000";
data_b(397) <= "0000000000";
data_b(398) <= "0000000000";
data_b(399) <= "0000000000";
----------------------------------25
data_b(400) <= "0000000100";
data_b(401) <= "0000000000";
data_b(402) <= "0000000000";
data_b(403) <= "0000000000";
data_b(404) <= "0000000000";
data_b(405) <= "0000000000";
data_b(406) <= "0000000000";
data_b(407) <= "0000000000";
data_b(408) <= "0000000000";
data_b(409) <= "0000000000";
data_b(410) <= "0000000000";
data_b(411) <= "0000000000";
data_b(412) <= "0000000000";
data_b(413) <= "0000000000";
data_b(414) <= "0000000000";
data_b(415) <= "0000000000";
---------------------------------26
data_b(416) <= "0000000010";
data_b(417) <= "0000000000";
data_b(418) <= "0000000010";
data_b(419) <= "0000000000";
data_b(420) <= "0000000000";
data_b(421) <= "0000000000";
data_b(422) <= "0000000010";
data_b(423) <= "0000000000";
data_b(424) <= "0000000000";
data_b(425) <= "0000000000";
data_b(426) <= "0000000010";
data_b(427) <= "0000000000";
data_b(428) <= "0000000001";
data_b(429) <= "0000000000";
data_b(430) <= "0000000000";
data_b(431) <= "0000000000";
---------------------------------27
data_b(432) <= "0000000001";
data_b(433) <= "0000000000";
data_b(434) <= "0000000010";
data_b(435) <= "0000000000";
data_b(436) <= "0000000000";
data_b(437) <= "0000000000";
data_b(438) <= "0000000100";
data_b(439) <= "0000000000";
data_b(440) <= "0010000000";
data_b(441) <= "0010000000";
data_b(442) <= "0010000000";
data_b(443) <= "0010000000";
data_b(444) <= "0000000000";
data_b(445) <= "0000000000";
data_b(446) <= "0000000000";
data_b(447) <= "0000000000";
------------------------------28
data_b(448) <= "0000000100";
data_b(449) <= "0000000000";
data_b(450) <= "0000000100";
data_b(451) <= "0000000000";
data_b(452) <= "0000000000";
data_b(453) <= "0000000000";
data_b(454) <= "0000000100";
data_b(455) <= "0000000000";
data_b(456) <= "0000000000";
data_b(457) <= "0000000000";
data_b(458) <= "0000000100";
data_b(459) <= "0000000000";
data_b(460) <= "0000000010";
data_b(461) <= "0000000000";
data_b(462) <= "0000000001";
data_b(463) <= "0000000000";
------------------------------29
data_b(464) <= "0000000000";
data_b(465) <= "0000000000";
data_b(466) <= "0000000000";
data_b(467) <= "0000000000";
data_b(468) <= "0000000000";
data_b(469) <= "0000000000";
data_b(470) <= "0000000000";
data_b(471) <= "0000000000";
data_b(472) <= "0000000000";
data_b(473) <= "0000000000";
data_b(474) <= "0000000000";
data_b(475) <= "0000000000";
data_b(476) <= "0000000000";
data_b(477) <= "0000000000";
data_b(478) <= "0000000000";
data_b(479) <= "0000000000";
--------------------------------30
data_b(480) <= "0000000010";
data_b(481) <= "0000000000";
data_b(482) <= "0000000010";
data_b(483) <= "0000000000";
data_b(484) <= "0000000000";
data_b(485) <= "0000000000";
data_b(486) <= "0000000010";
data_b(487) <= "0000000000";
data_b(488) <= "0000000000";
data_b(489) <= "0000000000";
data_b(490) <= "0000000010";
data_b(491) <= "0000000000";
data_b(492) <= "0000000001";
data_b(493) <= "0000000000";
data_b(494) <= "0000000000";
data_b(495) <= "0000000000";
----------------------------------31
data_b(496) <= "0010000000";
data_b(497) <= "0000000000";
data_b(498) <= "0000000010";
data_b(499) <= "0000000000";
data_b(500) <= "0000000000";
data_b(501) <= "0000000000";
data_b(502) <= "0000000100";
data_b(503) <= "0000000000";
data_b(504) <= "0010000000";
data_b(505) <= "0010000000";
data_b(506) <= "0010000000";
data_b(507) <= "0010000000";
data_b(508) <= "0000000000";
data_b(509) <= "0000000000";
data_b(510) <= "0000000000";
data_b(511) <= "0000000000";
----------------------------------32
data_b(512) <= "1000000000";
data_b(513) <= "0000000000";
data_b(514) <= "1000000000";
data_b(515) <= "0000000000";
data_b(516) <= "0000000000";
data_b(517) <= "0000000000";
data_b(518) <= "1000000000";
data_b(519) <= "0000000000";
data_b(520) <= "0000000000";
data_b(521) <= "0000000000";
data_b(522) <= "1000000000";
data_b(523) <= "0000000000";
data_b(524) <= "1000000000";
data_b(525) <= "0000000000";
data_b(526) <= "0000000000";
data_b(527) <= "0000000000";
-----------------------------------33
data_b(528) <= "0000000001";
data_b(529) <= "0000000000";
data_b(530) <= "0000000000";
data_b(531) <= "0000000000";
data_b(532) <= "0000000000";
data_b(533) <= "0000000000";
data_b(534) <= "0000000000";
data_b(535) <= "0000000000";
data_b(536) <= "0010000000";
data_b(537) <= "0000000000";
data_b(538) <= "0000000000";
data_b(539) <= "0000000000";
data_b(540) <= "0000000000";
data_b(541) <= "0000000000";
data_b(542) <= "0000000000";
data_b(543) <= "0000000000";
---------------------------------34
data_b(544) <= "0000000100";
data_b(545) <= "0000000000";
data_b(546) <= "0000000000";
data_b(547) <= "0000000000";
data_b(548) <= "0000000000";
data_b(549) <= "0000000000";
data_b(550) <= "0010000000";
data_b(551) <= "0000000000";
data_b(552) <= "0000000000";
data_b(553) <= "0000000000";
data_b(554) <= "0000000000";
data_b(555) <= "0000000000";
data_b(556) <= "1000000000";
data_b(557) <= "0000000000";
data_b(558) <= "0000000000";
data_b(559) <= "0000000000";
----------------------------------35
data_b(560) <= "0000000000";
data_b(561) <= "0000000000";
data_b(562) <= "0100000000";
data_b(563) <= "0000000000";
data_b(564) <= "0000000000";
data_b(565) <= "0000000000";
data_b(566) <= "0010000000";
data_b(567) <= "0000000000";
data_b(568) <= "0000000000";
data_b(569) <= "0000000000";
data_b(570) <= "0010000000";
data_b(571) <= "0000000000";
data_b(572) <= "0100000000";
data_b(573) <= "0000000000";
data_b(574) <= "0000000000";
data_b(575) <= "0000000000";
----------------------------------36
data_b(576) <= "1000000000";
data_b(577) <= "0000000000";
data_b(578) <= "0000000000";
data_b(579) <= "0100000000";
data_b(580) <= "0000000000";
data_b(581) <= "0000000000";
data_b(582) <= "0010000000";
data_b(583) <= "0000000000";
data_b(584) <= "0000000100";
data_b(585) <= "0000000000";
data_b(586) <= "0000000000";
data_b(587) <= "0000000000";
data_b(588) <= "0010000000";
data_b(589) <= "0000000000";
data_b(590) <= "0000000100";
data_b(591) <= "0000000000";
-----------------------------------37
data_b(592) <= "0000000000";
data_b(593) <= "0000000000";
data_b(594) <= "0000000100";
data_b(595) <= "0000000000";
data_b(596) <= "0000000000";
data_b(597) <= "0000000000";
data_b(598) <= "0100000000";
data_b(599) <= "0000000000";
data_b(600) <= "0010000000";
data_b(601) <= "0000000000";
data_b(602) <= "1000000000";
data_b(603) <= "0000000000";
data_b(604) <= "0000000000";
data_b(605) <= "0000000000";
data_b(606) <= "0000000000";
data_b(607) <= "0000000000";
-----------------------------------38
data_b(608) <= "0000000100";
data_b(609) <= "0000000000";
data_b(610) <= "0000000000";
data_b(611) <= "0000000000";
data_b(612) <= "0000000000";
data_b(613) <= "0000000000";
data_b(614) <= "0010000000";
data_b(615) <= "0000000000";
data_b(616) <= "0000000000";
data_b(617) <= "0000000000";
data_b(618) <= "0000000000";
data_b(619) <= "0000000000";
data_b(620) <= "1000000000";
data_b(621) <= "0000000000";
data_b(622) <= "0000000000";
data_b(623) <= "0000000000";
----------------------------------39
data_b(624) <= "0000000000";
data_b(625) <= "0000000000";
data_b(626) <= "0000000100";
data_b(627) <= "0000000000";
data_b(628) <= "0000000000";
data_b(629) <= "0000000000";
data_b(630) <= "0000000010";
data_b(631) <= "0000000000";
data_b(632) <= "0000000000";
data_b(633) <= "0000000000";
data_b(634) <= "0000000010";
data_b(635) <= "0000000000";
data_b(636) <= "0000000100";
data_b(637) <= "0000000000";
data_b(638) <= "0000000000";
data_b(639) <= "0000000000";
-----------------------------------40
data_b(640) <= "0010000000";
data_b(641) <= "0000000000";
data_b(642) <= "0000000000";
data_b(643) <= "0000000100";
data_b(644) <= "0000000000";
data_b(645) <= "0000000000";
data_b(646) <= "0000000010";
data_b(647) <= "0000000000";
data_b(648) <= "0000000001";
data_b(649) <= "0000000000";
data_b(650) <= "0000000000";
data_b(651) <= "0000000000";
data_b(652) <= "0000000010";
data_b(653) <= "0000000000";
data_b(654) <= "0000000001";
data_b(655) <= "0000000000";
---------------------------------41
data_b(656) <= "0000000000";
data_b(657) <= "0000000000";
data_b(658) <= "0000000001";
data_b(659) <= "0000000000";
data_b(660) <= "0000000000";
data_b(661) <= "0000000000";
data_b(662) <= "0000000100";
data_b(663) <= "0000000000";
data_b(664) <= "0000000010";
data_b(665) <= "0000000000";
data_b(666) <= "0010000000";
data_b(667) <= "0000000000";
data_b(668) <= "0000000000";
data_b(669) <= "0000000000";
data_b(670) <= "0000000000";
data_b(671) <= "0000000000";
-----------------------------------42
data_b(672) <= "0000000001";
data_b(673) <= "0000000000";
data_b(674) <= "0000000010";
data_b(675) <= "0000000000";
data_b(676) <= "0000000000";
data_b(677) <= "0000000000";
data_b(678) <= "0010000000";
data_b(679) <= "0000000000";
data_b(680) <= "0000000000";
data_b(681) <= "0000000000";
data_b(682) <= "0000000000";
data_b(683) <= "0000000000";
data_b(684) <= "0010000000";
data_b(685) <= "0000000000";
data_b(686) <= "0000000000";
data_b(687) <= "0000000000";
------------------------------------43
data_b(688) <= "0010000000";
data_b(689) <= "0000000000";
data_b(690) <= "0000000001";
data_b(691) <= "0000000000";
data_b(692) <= "0000000000";
data_b(693) <= "0000000000";
data_b(694) <= "0000000001";
data_b(695) <= "0000000000";
data_b(696) <= "0010000000";
data_b(697) <= "0000000000";
data_b(698) <= "0000000000";
data_b(699) <= "0000000000";
data_b(700) <= "0000000000";
data_b(701) <= "0000000000";
data_b(702) <= "0000000000";
data_b(703) <= "0000000000";
--------------------------------44
data_b(704) <= "0010000000";
data_b(705) <= "0000000000";
data_b(706) <= "0000000000";
data_b(707) <= "0000000001";
data_b(708) <= "0000000000";
data_b(709) <= "0000000000";
data_b(710) <= "0000000001";
data_b(711) <= "0000000000";
data_b(712) <= "0000000001";
data_b(713) <= "0000000000";
data_b(714) <= "0000000000";
data_b(715) <= "0000000010";
data_b(716) <= "0000000000";
data_b(717) <= "0000000000";
data_b(718) <= "0000000100";
data_b(719) <= "0000000000";
-------------------------------45
data_b(720) <= "0000000001";
data_b(721) <= "0000000000";
data_b(722) <= "0000000010";
data_b(723) <= "0000000000";
data_b(724) <= "0000000000";
data_b(725) <= "0000000000";
data_b(726) <= "0000000100";
data_b(727) <= "0000000000";
data_b(728) <= "0010000000";
data_b(729) <= "0000000000";
data_b(730) <= "0000000000";
data_b(731) <= "0000000000";
data_b(732) <= "0000000000";
data_b(733) <= "0000000000";
data_b(734) <= "0000000000";
data_b(735) <= "0000000000";
-------------------------------46
data_b(736) <= "0000000001";
data_b(737) <= "0000000000";
data_b(738) <= "0000000010";
data_b(739) <= "0000000000";
data_b(740) <= "0000000000";
data_b(741) <= "0000000000";
data_b(742) <= "0000000100";
data_b(743) <= "0000000000";
data_b(744) <= "0000000000";
data_b(745) <= "0000000000";
data_b(746) <= "0000000000";
data_b(747) <= "0000000000";
data_b(748) <= "0000000100";
data_b(749) <= "0000000000";
data_b(750) <= "0000000000";
data_b(751) <= "0000000000";
----------------------------47
data_b(752) <= "0010000000";
data_b(753) <= "0000000000";
data_b(754) <= "0000000001";
data_b(755) <= "0000000000";
data_b(756) <= "0000000000";
data_b(757) <= "0000000000";
data_b(758) <= "0000000001";
data_b(759) <= "0000000000";
data_b(760) <= "0010000000";
data_b(761) <= "0000000000";
data_b(762) <= "0000000000";
data_b(763) <= "0000000000";
data_b(764) <= "0000000000";
data_b(765) <= "0000000000";
data_b(766) <= "0000000000";
data_b(767) <= "0000000000";
--------------------------------48
data_b(768) <= "0010000000";
data_b(769) <= "0000000000";
data_b(770) <= "0000000001";
data_b(771) <= "0000000000";
data_b(772) <= "0000000000";
data_b(773) <= "0000000000";
data_b(774) <= "0000000001";
data_b(775) <= "0000000000";
data_b(776) <= "0000000001";
data_b(777) <= "0000000000";
data_b(778) <= "0000000000";
data_b(779) <= "0000000010";
data_b(780) <= "0000000000";
data_b(781) <= "0000000000";
data_b(782) <= "0000000100";
data_b(783) <= "0000000000";
-------------------------------49
data_b(784) <= "0000000010";
data_b(785) <= "0000000000";
data_b(786) <= "0000000000";
data_b(787) <= "0000000000";
data_b(788) <= "0000000000";
data_b(789) <= "0000000000";
data_b(790) <= "0000000000";
data_b(791) <= "0000000000";
data_b(792) <= "0000000000";
data_b(793) <= "0000000000";
data_b(794) <= "0000000000";
data_b(795) <= "0000000000";
data_b(796) <= "0000000000";
data_b(797) <= "0000000000";
data_b(798) <= "0000000000";
data_b(799) <= "0000000000";
----------------------------50
data_b(800) <= "0000000001";
data_b(801) <= "0000000000";
data_b(802) <= "0000000010";
data_b(803) <= "0000000000";
data_b(804) <= "0000000000";
data_b(805) <= "0000000000";
data_b(806) <= "0010000000";
data_b(807) <= "0000000000";
data_b(808) <= "0000000000";
data_b(809) <= "0000000000";
data_b(810) <= "0000000000";
data_b(811) <= "0000000000";
data_b(812) <= "0010000000";
data_b(813) <= "0000000000";
data_b(814) <= "0000000000";
data_b(815) <= "0000000000";
----------------------------------51
data_b(816) <= "0010000000";
data_b(817) <= "0000000000";
data_b(818) <= "0000000001";
data_b(819) <= "0000000000";
data_b(820) <= "0000000000";
data_b(821) <= "0000000000";
data_b(822) <= "0000000001";
data_b(823) <= "0000000000";
data_b(824) <= "0010000000";
data_b(825) <= "0000000000";
data_b(826) <= "0000000000";
data_b(827) <= "0000000000";
data_b(828) <= "0000000000";
data_b(829) <= "0000000000";
data_b(830) <= "0000000000";
data_b(831) <= "0000000000";
--------------------------------52
data_b(832) <= "0010000000";
data_b(833) <= "0000000000";
data_b(834) <= "0000000000";
data_b(835) <= "0000000001";
data_b(836) <= "0000000000";
data_b(837) <= "0000000000";
data_b(838) <= "0000000001";
data_b(839) <= "0000000000";
data_b(840) <= "0000000001";
data_b(841) <= "0000000000";
data_b(842) <= "0000000000";
data_b(843) <= "0000000010";
data_b(844) <= "0000000000";
data_b(845) <= "0000000000";
data_b(846) <= "0000000100";
data_b(847) <= "0000000000";
------------------------------53
data_b(848) <= "0000000001";
data_b(849) <= "0000000000";
data_b(850) <= "0000000010";
data_b(851) <= "0000000000";
data_b(852) <= "0000000000";
data_b(853) <= "0000000000";
data_b(854) <= "0000000100";
data_b(855) <= "0000000000";
data_b(856) <= "0010000000";
data_b(857) <= "0000000000";
data_b(858) <= "0000000000";
data_b(859) <= "0000000000";
data_b(860) <= "0000000000";
data_b(861) <= "0000000000";
data_b(862) <= "0000000000";
data_b(863) <= "0000000000";
------------------------------54
data_b(864) <= "0000000001";
data_b(865) <= "0000000000";
data_b(866) <= "0000000010";
data_b(867) <= "0000000000";
data_b(868) <= "0000000000";
data_b(869) <= "0000000000";
data_b(870) <= "0010000000";
data_b(871) <= "0000000000";
data_b(872) <= "0000000000";
data_b(873) <= "0000000000";
data_b(874) <= "0000000000";
data_b(875) <= "0000000000";
data_b(876) <= "0010000000";
data_b(877) <= "0000000000";
data_b(878) <= "0000000000";
data_b(879) <= "0000000000";
-----------------------------55
data_b(880) <= "0010000000";
data_b(881) <= "0000000000";
data_b(882) <= "0000000001";
data_b(883) <= "0000000000";
data_b(884) <= "0000000000";
data_b(885) <= "0000000000";
data_b(886) <= "0000000001";
data_b(887) <= "0000000000";
data_b(888) <= "0010000000";
data_b(889) <= "0000000000";
data_b(890) <= "0000000000";
data_b(891) <= "0000000000";
data_b(892) <= "0000000000";
data_b(893) <= "0000000000";
data_b(894) <= "0000000000";
data_b(895) <= "0000000000";
--------------------------------56
data_b(896) <= "0010000000";
data_b(897) <= "0000000000";
data_b(898) <= "0000000001";
data_b(899) <= "0000000000";
data_b(900) <= "0000000000";
data_b(901) <= "0000000000";
data_b(902) <= "0000000001";
data_b(903) <= "0000000000";
data_b(904) <= "0000000001";
data_b(905) <= "0000000000";
data_b(906) <= "0000000000";
data_b(907) <= "0000000010";
data_b(908) <= "0000000000";
data_b(909) <= "0000000000";
data_b(910) <= "0000000100";
data_b(911) <= "0000000000";
-------------------------------57
data_b(912) <= "0000000100";
data_b(913) <= "0000000000";
data_b(914) <= "0000000000";
data_b(915) <= "0000000000";
data_b(916) <= "0000000000";
data_b(917) <= "0000000000";
data_b(918) <= "0000000000";
data_b(919) <= "0000000000";
data_b(920) <= "0000000000";
data_b(921) <= "0000000000";
data_b(922) <= "0000000000";
data_b(923) <= "0000000000";
data_b(924) <= "0000000000";
data_b(925) <= "0000000000";
data_b(926) <= "0000000000";
data_b(927) <= "0000000000";
-----------------------------58
data_b(928) <= "0000000100";
data_b(939) <= "0000000000";
data_b(930) <= "0000000100";
data_b(931) <= "0000000000";
data_b(932) <= "0000000000";
data_b(933) <= "0000000000";
data_b(934) <= "0000000100";
data_b(935) <= "0000000000";
data_b(936) <= "0000000000";
data_b(937) <= "0000000000";
data_b(938) <= "0000000100";
data_b(939) <= "0000000000";
data_b(940) <= "0000000010";
data_b(941) <= "0000000000";
data_b(942) <= "0000000000";
data_b(943) <= "0000000000";
-------------------------------59
data_b(944) <= "0000000001";
data_b(945) <= "0000000000";
data_b(946) <= "0000000010";
data_b(947) <= "0000000000";
data_b(948) <= "0000000000";
data_b(949) <= "0000000000";
data_b(950) <= "0000000100";
data_b(951) <= "0000000000";
data_b(952) <= "0010000000";
data_b(953) <= "0010000000";
data_b(954) <= "0010000000";
data_b(955) <= "0010000000";
data_b(956) <= "0000000000";
data_b(957) <= "0000000000";
data_b(958) <= "0000000000";
data_b(959) <= "0000000000";
-----------------------------60
data_b(960) <= "0000000100";
data_b(961) <= "0000000000";
data_b(962) <= "0000000100";
data_b(963) <= "0000000000";
data_b(964) <= "0000000000";
data_b(965) <= "0000000000";
data_b(966) <= "0000000100";
data_b(967) <= "0000000000";
data_b(968) <= "0000000000";
data_b(969) <= "0000000000";
data_b(970) <= "0000000100";
data_b(971) <= "0000000000";
data_b(972) <= "0000000010";
data_b(973) <= "0000000000";
data_b(974) <= "0000000001";
data_b(975) <= "0000000000";
-------------------------------61
data_b(976) <= "0000000000";
data_b(977) <= "0000000000";
data_b(978) <= "0000000000";
data_b(979) <= "0000000000";
data_b(980) <= "0000000100";
data_b(981) <= "0000000000";
data_b(982) <= "0000000010";
data_b(983) <= "0000000000";
data_b(984) <= "0010000000";
data_b(985) <= "0000000000";
data_b(986) <= "0000000010";
data_b(987) <= "0000000000";
data_b(988) <= "0000000001";
data_b(989) <= "0000000000";
data_b(990) <= "0010000000";
data_b(991) <= "0000000000";
----------------------------62
data_b(992) <= "0000000010";
data_b(993) <= "0000000000";
data_b(994) <= "0000000010";
data_b(995) <= "0000000000";
data_b(996) <= "0000000000";
data_b(997) <= "0000000000";
data_b(998) <= "0000000010";
data_b(999) <= "0000000000";
data_b(1000) <= "0000000000";
data_b(1001) <= "0000000000";
data_b(1002) <= "0000000010";
data_b(1003) <= "0000000000";
data_b(1004) <= "0000000001";
data_b(1005) <= "0000000000";
data_b(1006) <= "0000000000";
data_b(1007) <= "0000000000";
---------------------------------63
data_b(1008) <= "0000000001";
data_b(1009) <= "0000000000";
data_b(1010) <= "0000000010";
data_b(1011) <= "0000000000";
data_b(1012) <= "0000000000";
data_b(1013) <= "0000000000";
data_b(1014) <= "0000000100";
data_b(1015) <= "0000000000";
data_b(1016) <= "0010000000";
data_b(1017) <= "0010000000";
data_b(1018) <= "0010000000";
data_b(1019) <= "0010000000";
data_b(1020) <= "0000000000";
data_b(1021) <= "0000000000";
data_b(1022) <= "0000000000";
data_b(1023) <= "0000000000";
-----------------------------64
data_b(1024) <= "0000000001";
data_b(1025) <= "0000000000";
data_b(1026) <= "0000000001";
data_b(1027) <= "0000000000";
data_b(1028) <= "0000000000";
data_b(1029) <= "0000000000";
data_b(1030) <= "0000000001";
data_b(1031) <= "0000000000";
data_b(1032) <= "0000000000";
data_b(1033) <= "0000000000";
data_b(1034) <= "0000000010";
data_b(1035) <= "0000000000";
data_b(1036) <= "0000000001";
data_b(1037) <= "0000000000";
data_b(1038) <= "0000000000";
data_b(1039) <= "0000000000";
--------------------------------65
data_b(1040) <= "0000000001";
data_b(1041) <= "0000000000";
data_b(1042) <= "0000000000";
data_b(1043) <= "0000000000";
data_b(1044) <= "0000000000";
data_b(1045) <= "0000000000";
data_b(1046) <= "0000000000";
data_b(1047) <= "0000000000";
data_b(1048) <= "0010000000";
data_b(1049) <= "0000000000";
data_b(1050) <= "0000000000";
data_b(1051) <= "0000000000";
data_b(1052) <= "0000000000";
data_b(1053) <= "0000000000";
data_b(1054) <= "0000000000";
data_b(1055) <= "0000000000";
--------------------------------66
data_b(1056) <= "0000000001";
data_b(1057) <= "0000000000";
data_b(1058) <= "0000000010";
data_b(1059) <= "0000000000";
data_b(1060) <= "0000000000";
data_b(1061) <= "0000000000";
data_b(1062) <= "0010000000";
data_b(1063) <= "0000000000";
data_b(1064) <= "0000000000";
data_b(1065) <= "0000000000";
data_b(1066) <= "0000000000";
data_b(1067) <= "0000000000";
data_b(1068) <= "0010000000";
data_b(1069) <= "0000000000";
data_b(1070) <= "0000000000";
data_b(1071) <= "0000000000";
------------------------------------67
data_b(1072) <= "0010000000";
data_b(1073) <= "0000000000";
data_b(1074) <= "0000000001";
data_b(1075) <= "0000000000";
data_b(1076) <= "0000000000";
data_b(1077) <= "0000000000";
data_b(1078) <= "0000000001";
data_b(1079) <= "0000000000";
data_b(1080) <= "0010000000";
data_b(1081) <= "0000000000";
data_b(1082) <= "0000000000";
data_b(1083) <= "0000000000";
data_b(1084) <= "0000000000";
data_b(1085) <= "0000000000";
data_b(1086) <= "0000000000";
data_b(1087) <= "0000000000";
----------------------------------68
data_b(1088) <= "0010000000";
data_b(1089) <= "0000000000";
data_b(1090) <= "0000000000";
data_b(1091) <= "0000000001";
data_b(1092) <= "0000000000";
data_b(1093) <= "0000000000";
data_b(1094) <= "0000000001";
data_b(1095) <= "0000000000";
data_b(1096) <= "0000000001";
data_b(1097) <= "0000000000";
data_b(1098) <= "0000000000";
data_b(1099) <= "0000000010";
data_b(1100) <= "0000000000";
data_b(1101) <= "0000000000";
data_b(1102) <= "0000000100";
data_b(1103) <= "0000000000";
------------------------------69
data_b(1104) <= "0000000001";
data_b(1105) <= "0000000000";
data_b(1106) <= "0000000010";
data_b(1107) <= "0000000000";
data_b(1108) <= "0000000000";
data_b(1109) <= "0000000000";
data_b(1110) <= "0000000100";
data_b(1111) <= "0000000000";
data_b(1112) <= "0010000000";
data_b(1113) <= "0000000000";
data_b(1114) <= "0000000000";
data_b(1115) <= "0000000000";
data_b(1116) <= "0000000000";
data_b(1117) <= "0000000000";
data_b(1118) <= "0000000000";
data_b(1119) <= "0000000000";
--------------------------------70
data_b(1120) <= "0000000001";
data_b(1121) <= "0000000000";
data_b(1122) <= "0000000010";
data_b(1123) <= "0000000000";
data_b(1124) <= "0000000000";
data_b(1125) <= "0000000000";
data_b(1126) <= "0010000000";
data_b(1127) <= "0000000000";
data_b(1128) <= "0000000000";
data_b(1129) <= "0000000000";
data_b(1130) <= "0000000000";
data_b(1131) <= "0000000000";
data_b(1132) <= "0010000000";
data_b(1133) <= "0000000000";
data_b(1134) <= "0000000000";
data_b(1135) <= "0000000000";
-----------------------------71
data_b(1136) <= "0010000000";
data_b(1137) <= "0000000000";
data_b(1138) <= "0000000001";
data_b(1139) <= "0000000000";
data_b(1140) <= "0000000000";
data_b(1141) <= "0000000000";
data_b(1142) <= "0000000001";
data_b(1143) <= "0000000000";
data_b(1144) <= "0010000000";
data_b(1145) <= "0000000000";
data_b(1146) <= "0000000000";
data_b(1147) <= "0000000000";
data_b(1148) <= "0000000000";
data_b(1149) <= "0000000000";
data_b(1150) <= "0000000000";
data_b(1151) <= "0000000000";
---------------------------------72
data_b(1152) <= "0010000000";
data_b(1153) <= "0000000000";
data_b(1154) <= "0000000001";
data_b(1155) <= "0000000000";
data_b(1156) <= "0000000000";
data_b(1157) <= "0000000000";
data_b(1158) <= "0000000001";
data_b(1159) <= "0000000000";
data_b(1160) <= "0000000001";
data_b(1161) <= "0000000000";
data_b(1162) <= "0000000000";
data_b(1163) <= "0000000010";
data_b(1164) <= "0000000000";
data_b(1165) <= "0000000000";
data_b(1166) <= "0000000100";
data_b(1167) <= "0000000000";
--------------------------------73
data_b(1168) <= "0000000100";
data_b(1169) <= "0000000000";
data_b(1170) <= "0000000000";
data_b(1171) <= "0000000000";
data_b(1172) <= "0000000000";
data_b(1173) <= "0000000000";
data_b(1174) <= "0000000000";
data_b(1175) <= "0000000000";
data_b(1176) <= "0000000000";
data_b(1177) <= "0000000000";
data_b(1178) <= "0000000000";
data_b(1179) <= "0000000000";
data_b(1180) <= "0000000000";
data_b(1181) <= "0000000000";
data_b(1182) <= "0000000000";
data_b(1183) <= "0000000000";
-------------------------------------74
data_b(1184) <= "0000000001";
data_b(1185) <= "0000000000";
data_b(1186) <= "0000000010";
data_b(1187) <= "0000000000";
data_b(1188) <= "0000000000";
data_b(1189) <= "0000000000";
data_b(1190) <= "0010000000";
data_b(1191) <= "0000000000";
data_b(1192) <= "0000000000";
data_b(1193) <= "0000000000";
data_b(1194) <= "0000000000";
data_b(1195) <= "0000000000";
data_b(1196) <= "0010000000";
data_b(1197) <= "0000000000";
data_b(1198) <= "0000000000";
data_b(1199) <= "0000000000";
-------------------------------------75
data_b(1200) <= "0010000000";
data_b(1201) <= "0000000000";
data_b(1202) <= "0000000001";
data_b(1203) <= "0000000000";
data_b(1204) <= "0000000000";
data_b(1205) <= "0000000000";
data_b(1206) <= "0000000001";
data_b(1207) <= "0000000000";
data_b(1208) <= "0010000000";
data_b(1209) <= "0000000000";
data_b(1210) <= "0000000000";
data_b(1211) <= "0000000000";
data_b(1212) <= "0000000000";
data_b(1213) <= "0000000000";
data_b(1214) <= "0000000000";
data_b(1215) <= "0000000000";
----------------------------------76
data_b(1216) <= "0010000000";
data_b(1217) <= "0000000000";
data_b(1218) <= "0000000000";
data_b(1219) <= "0000000001";
data_b(1220) <= "0000000000";
data_b(1221) <= "0000000000";
data_b(1222) <= "0000000001";
data_b(1223) <= "0000000000";
data_b(1224) <= "0000000001";
data_b(1225) <= "0000000000";
data_b(1226) <= "0000000000";
data_b(1227) <= "0000000010";
data_b(1228) <= "0000000000";
data_b(1229) <= "0000000000";
data_b(1230) <= "0000000100";
data_b(1231) <= "0000000000";
-------------------------------77
data_b(1232) <= "0000000001";
data_b(1233) <= "0000000000";
data_b(1234) <= "0000000010";
data_b(1235) <= "0000000000";
data_b(1236) <= "0000000000";
data_b(1237) <= "0000000000";
data_b(1238) <= "0000000100";
data_b(1239) <= "0000000000";
data_b(1240) <= "0010000000";
data_b(1241) <= "0000000000";
data_b(1242) <= "0000000000";
data_b(1243) <= "0000000000";
data_b(1244) <= "0000000000";
data_b(1245) <= "0000000000";
data_b(1246) <= "0000000000";
data_b(1247) <= "0000000000";
-------------------------------78
data_b(1248) <= "0000000001";
data_b(1249) <= "0000000000";
data_b(1250) <= "0000000010";
data_b(1251) <= "0000000000";
data_b(1252) <= "0000000000";
data_b(1253) <= "0000000000";
data_b(1254) <= "0010000000";
data_b(1255) <= "0000000000";
data_b(1256) <= "0000000000";
data_b(1257) <= "0000000000";
data_b(1258) <= "0000000000";
data_b(1259) <= "0000000000";
data_b(1260) <= "0010000000";
data_b(1261) <= "0000000000";
data_b(1262) <= "0000000000";
data_b(1263) <= "0000000000";
-----------------------------79
data_b(1264) <= "0010000000";
data_b(1265) <= "0000000000";
data_b(1266) <= "0000000001";
data_b(1267) <= "0000000000";
data_b(1268) <= "0000000000";
data_b(1269) <= "0000000000";
data_b(1270) <= "0000000001";
data_b(1271) <= "0000000000";
data_b(1272) <= "0001000000";
data_b(1273) <= "0000000000";
data_b(1274) <= "0000000000";
data_b(1275) <= "0000000000";
data_b(1276) <= "0000000000";
data_b(1277) <= "0000000000";
data_b(1278) <= "0000000000";
data_b(1279) <= "0000000000";
----------------------------------80
data_b(1280) <= "0001000000";
data_b(1281) <= "0000000000";
data_b(1282) <= "0000000001";
data_b(1283) <= "0000000000";
data_b(1284) <= "0000000000";
data_b(1285) <= "0000000000";
data_b(1286) <= "0000000001";
data_b(1287) <= "0000000000";
data_b(1288) <= "0000000001";
data_b(1289) <= "0000000000";
data_b(1290) <= "0000000000";
data_b(1291) <= "0000000010";
data_b(1292) <= "0000000000";
data_b(1293) <= "0000000000";
data_b(1294) <= "0000000100";
data_b(1295) <= "0000000000";
--------------------------------81
data_b(1296) <= "0000000010";
data_b(1297) <= "0000000000";
data_b(1298) <= "0000000000";
data_b(1299) <= "0000000000";
data_b(1300) <= "0000000000";
data_b(1301) <= "0000000000";
data_b(1302) <= "0000000000";
data_b(1303) <= "0000000000";
data_b(1304) <= "0000000000";
data_b(1305) <= "0000000000";
data_b(1306) <= "0000000000";
data_b(1307) <= "0000000000";
data_b(1308) <= "0000000000";
data_b(1309) <= "0000000000";
data_b(1310) <= "0000000000";
data_b(1311) <= "0000000000";
-----------------------------------82
data_b(1312) <= "0000000001";
data_b(1313) <= "0000000000";
data_b(1314) <= "0000000000";
data_b(1315) <= "0000000000";
data_b(1316) <= "0000000000";
data_b(1317) <= "0000000000";
data_b(1318) <= "0000000010";
data_b(1319) <= "0000000000";
data_b(1320) <= "0000000000";
data_b(1321) <= "0000000000";
data_b(1322) <= "0000000000";
data_b(1323) <= "0000000000";
data_b(1324) <= "0000000100";
data_b(1325) <= "0000000000";
data_b(1326) <= "0000000000";
data_b(1327) <= "0000000000";
------------------------------83
data_b(1328) <= "0000000100";
data_b(1329) <= "0000000000";
data_b(1330) <= "0000000000";
data_b(1331) <= "0000000010";
data_b(1332) <= "0000000000";
data_b(1333) <= "0000000000";
data_b(1334) <= "0000000100";
data_b(1335) <= "0000000000";
data_b(1336) <= "0000000100";
data_b(1337) <= "0000000000";
data_b(1338) <= "0000000000";
data_b(1339) <= "0000000010";
data_b(1340) <= "0000000000";
data_b(1341) <= "0000000000";
data_b(1342) <= "0000000100";
data_b(1343) <= "0000000000";
------------------------------84
data_b(1344) <= "0000000010";
data_b(1345) <= "0000000010";
data_b(1346) <= "0000000010";
data_b(1347) <= "0000000010";
data_b(1348) <= "0000000000";
data_b(1349) <= "0000000000";
data_b(1350) <= "0000000000";
data_b(1351) <= "0000000000";
data_b(1352) <= "0000000100";
data_b(1353) <= "0000000100";
data_b(1354) <= "0000000100";
data_b(1355) <= "0000000100";
data_b(1356) <= "0000000000";
data_b(1357) <= "0000000000";
data_b(1358) <= "0000000000";
data_b(1359) <= "0000000000";
-----------------------------------85


----------------------------
--------------------1
scale2(15) <= d_3;
scale2(16) <=  r;
scale2(17) <=  d_3;
scale2(18) <=  d_3;
scale2(19) <=  r;
scale2(20) <=  r;
scale2(21) <=  d_3;
scale2(22) <=  d_3;
scale2(23) <=  r;
scale2(24) <=  r;
scale2(25) <=  d_3;
scale2(26) <=  r;
scale2(27) <=  d_3;
scale2(28) <=  d_3;
scale2(29) <=  d_3;
scale2(30) <=  r;
--------------------2
scale2(31) <= g_3;
scale2(32) <= g_3;
scale2(33) <= g_3;
scale2(34) <= g_3;
scale2(35) <= r;
scale2(36) <= r;
scale2(37) <= r;
scale2(38) <= r;
scale2(39) <= g_2;
scale2(40) <= g_2;
scale2(41) <= g_2;
scale2(42) <= g_2;
scale2(43) <= r;
scale2(44) <= r;
scale2(45) <= r;
scale2(46) <= r;
--------------------3
scale2(47) <= g_3;
scale2(48) <= g_3;
scale2(49) <= g_3;
scale2(50) <= g_3;
scale2(51) <= r;
scale2(52) <= r;
scale2(53) <= e_3;
scale2(54) <= e_3;
scale2(55) <= e_3;
scale2(56) <= e_3;
scale2(57) <= r;
scale2(58) <= r;
scale2(59) <= c_3;
scale2(60) <= c_3;
scale2(61) <= c_3;
scale2(62) <= c_3;
--------------------4
scale2(63) <= r;
scale2(64) <= r;
scale2(65) <= f_3;
scale2(66) <= f_3;
scale2(67) <= f_3;
scale2(68) <= r;
scale2(69) <= g_3;
scale2(70) <= g_3;
scale2(71) <= g_3;
scale2(72) <= r;
scale2(73) <= gm_3;
scale2(74) <= r;
scale2(75) <= f_3;
scale2(76) <= f_3;
scale2(77) <= f_3;
scale2(78) <= r;
--------------------5
scale2(79) <= e_3;
scale2(80) <= e_3;
scale2(81) <= r;
scale2(82) <= c_4;
scale2(83) <= c_4;
scale2(84) <= r;
scale2(85) <= e_4;
scale2(86) <= r;
scale2(87) <= f_4;
scale2(88) <= f_4;
scale2(89) <= f_4;
scale2(90) <= r;
scale2(91) <= d_4;
scale2(92) <= r;
scale2(93) <= e_4;
scale2(94) <= e_4;
-------------------6
scale2(95) <= r;
scale2(96) <= r;
scale2(97) <= c_4;
scale2(98) <= c_4;
scale2(99) <= c_4;
scale2(100) <= r;
scale2(101) <= a_4;
scale2(102) <= r;
scale2(103) <= b_4;
scale2(104) <= r;
scale2(105) <= g_4;
scale2(106) <= g_4;
scale2(107) <= g_4;
scale2(108) <= g_4;
scale2(109) <= r;
scale2(110) <= r;
--------------------7
scale2(111) <= g_3;
scale2(112) <= g_3;
scale2(113) <= g_3;
scale2(114) <= g_3;
scale2(115) <= r;
scale2(116) <= r;
scale2(117) <= e_3;
scale2(118) <= e_3;
scale2(119) <= e_3;
scale2(120) <= e_3;
scale2(121) <= r;
scale2(122) <= r;
scale2(123) <= c_3;
scale2(124) <= c_3;
scale2(125) <= c_3;
scale2(126) <= c_3;
--------------------8
scale2(127) <= r;
scale2(128) <= r;
scale2(129) <= f_3;
scale2(130) <= f_3;
scale2(131) <= f_3;
scale2(132) <= r;
scale2(133) <= g_3;
scale2(134) <= g_3;
scale2(135) <= g_3;
scale2(136) <= r;
scale2(137) <= gm_3;
scale2(138) <= r;
scale2(139) <= f_3;
scale2(140) <= f_3;
scale2(141) <= f_3;
scale2(142) <= r;
--------------------9
scale2(143) <= e_3;
scale2(144) <= e_3;
scale2(145) <= r;
scale2(146) <= c_4;
scale2(147) <= c_4;
scale2(148) <= r;
scale2(149) <= e_4;
scale2(150) <= r;
scale2(151) <= f_4;
scale2(152) <= f_4;
scale2(153) <= f_4;
scale2(154) <= r;
scale2(155) <= d_4;
scale2(156) <= r;
scale2(157) <= e_4;
scale2(158) <= e_4;
--------------------10
scale2(159) <= r;
scale2(160) <= r;
scale2(161) <= c_4;
scale2(162) <= c_4;
scale2(163) <= c_4;
scale2(164) <= r;
scale2(165) <= a_4;
scale2(166) <= r;
scale2(167) <= b_4;
scale2(168) <= r;
scale2(169) <= g_4;
scale2(170) <= g_4;
scale2(171) <= g_4;
scale2(172) <= g_4;
scale2(173) <= r;
scale2(174) <= r;
--------------------11
scale2(175) <= c_3;
scale2(176) <= c_3;
scale2(177) <= c_3;
scale2(178) <= c_3;
scale2(179) <= r;
scale2(180) <= r;
scale2(181) <= g_3;
scale2(182) <= g_3;
scale2(183) <= r;
scale2(184) <= r;
scale2(185) <= r;
scale2(186) <= r;
scale2(187) <= c_4;
scale2(188) <= c_4;
scale2(189) <= c_4;
scale2(190) <= r;
--------------------12
scale2(191) <= f_3;
scale2(192) <= f_3;
scale2(193) <= f_3;
scale2(194) <= f_3;
scale2(195) <= r;
scale2(196) <= r;
scale2(197) <= c_4;
scale2(198) <= r;
scale2(199) <= c_4;
scale2(200) <= c_4;
scale2(201) <= c_4;
scale2(202) <= r;
scale2(203) <= f_3;
scale2(204) <= f_3;
scale2(205) <= f_3;
scale2(206) <= r;
--------------------13
scale2(207) <= c_3;
scale2(208) <= c_3;
scale2(209) <= c_3;
scale2(210) <= c_3;
scale2(211) <= r;
scale2(212) <= r;
scale2(213) <= e_3;
scale2(214) <= e_3;
scale2(215) <= r;
scale2(216) <= r;
scale2(217) <= r;
scale2(218) <= r;
scale2(219) <= g_3;
scale2(220) <= r;
scale2(221) <= c_4;
scale2(222) <= c_4;
--------------------14
scale2(223) <= r;
scale2(224) <= r;
scale2(225) <= r;
scale2(226) <= r;
scale2(227) <= r;
scale2(228) <= r;
scale2(229) <= r;
scale2(230) <= r;
scale2(231) <= r;
scale2(232) <= r;
scale2(233) <= r;
scale2(234) <= r;
scale2(235) <= g_3;
scale2(236) <= g_3;
scale2(237) <= g_3;
scale2(238) <= r;
--------------------15
scale2(239) <= c_3;
scale2(240) <= c_3;
scale2(241) <= c_3;
scale2(242) <= c_3;
scale2(243) <= r;
scale2(244) <= r;
scale2(245) <= g_3;
scale2(246) <= g_3;
scale2(247) <= r;
scale2(248) <= r;
scale2(249) <= r;
scale2(250) <= r;
scale2(251) <= c_4;
scale2(252) <= c_4;
scale2(253) <= c_4;
scale2(254) <= r;
--------------------16
scale2(255) <= f_3;
scale2(256) <= f_3;
scale2(257) <= f_3;
scale2(258) <= f_3;
scale2(259) <= r;
scale2(260) <= r;
scale2(261) <= c_4;
scale2(262) <= r;
scale2(263) <= c_4;
scale2(264) <= c_4;
scale2(265) <= c_4;
scale2(266) <= r;
scale2(267) <= f_3;
scale2(268) <= f_3;
scale2(269) <= f_3;
scale2(270) <= r;
--------------------17
scale2(271) <= c_3;
scale2(272) <= c_3;
scale2(273) <= c_3;
scale2(274) <= r;
scale2(275) <= am_3;
scale2(276) <= am_3;
scale2(277) <= am_3;
scale2(278) <= am_3;
scale2(279) <= r;
scale2(280) <= r;
scale2(281) <= am_4;
scale2(282) <= am_4;
scale2(283) <= am_4;
scale2(284) <= am_4;
scale2(285) <= r;
scale2(286) <= r;
--------------------18
scale2(287) <= c_4;
scale2(288) <= c_4;
scale2(289) <= c_4;
scale2(290) <= c_4;
scale2(291) <= r;
scale2(292) <= r;
scale2(293) <= g_3;
scale2(294) <= r;
scale2(295) <= g_3;
scale2(296) <= g_3;
scale2(297) <= g_3;
scale2(298) <= r;
scale2(299) <= c_3;
scale2(300) <= c_3;
scale2(301) <= c_3;
scale2(302) <= r;
--------------------19
scale2(303) <= c_3;
scale2(304) <= c_3;
scale2(305) <= c_3;
scale2(306) <= c_3;
scale2(307) <= r;
scale2(308) <= r;
scale2(309) <= g_3;
scale2(310) <= g_3;
scale2(311) <= r;
scale2(312) <= r;
scale2(313) <= r;
scale2(314) <= r;
scale2(315) <= c_4;
scale2(316) <= c_4;
scale2(317) <= c_4;
scale2(318) <= r;
--------------------20
scale2(319) <= f_3;
scale2(320) <= f_3;
scale2(321) <= f_3;
scale2(322) <= f_3;
scale2(323) <= r;
scale2(324) <= r;
scale2(325) <= c_4;
scale2(326) <= r;
scale2(327) <= c_4;
scale2(328) <= c_4;
scale2(329) <= c_4;
scale2(330) <= r;
scale2(331) <= f_3;
scale2(332) <= f_3;
scale2(333) <= f_3;
scale2(334) <= r;
--------------------21
scale2(335) <= c_3;
scale2(336) <= c_3;
scale2(337) <= c_3;
scale2(338) <= c_3;
scale2(339) <= r;
scale2(340) <= r;
scale2(341) <= e_3;
scale2(342) <= e_3;
scale2(343) <= r;
scale2(344) <= r;
scale2(345) <= r;
scale2(346) <= r;
scale2(347) <= g_3;
scale2(348) <= r;
scale2(349) <= c_4;
scale2(350) <= c_4;
--------------------22
scale2(351) <= r;
scale2(352) <= r;
scale2(353) <= r;
scale2(354) <= r;
scale2(355) <= r;
scale2(356) <= r;
scale2(357) <= r;
scale2(358) <= r;
scale2(359) <= r;
scale2(360) <= r;
scale2(361) <= r;
scale2(362) <= r;
scale2(363) <= g_3;
scale2(364) <= g_3;
scale2(365) <= g_3;
scale2(366) <= r;
--------------------23
scale2(367) <= c_3;
scale2(368) <= c_3;
scale2(369) <= c_3;
scale2(370) <= c_3;
scale2(371) <= r;
scale2(372) <= r;
scale2(373) <= g_3;
scale2(374) <= g_3;
scale2(375) <= r;
scale2(376) <= r;
scale2(377) <= r;
scale2(378) <= r;
scale2(379) <= c_4;
scale2(380) <= c_4;
scale2(381) <= c_4;
scale2(382) <= r;
--------------------24
scale2(383) <= f_3;
scale2(384) <= f_3;
scale2(385) <= f_3;
scale2(386) <= f_3;
scale2(387) <= r;
scale2(388) <= r;
scale2(389) <= c_4;
scale2(390) <= r;
scale2(391) <= c_4;
scale2(392) <= c_4;
scale2(393) <= c_4;
scale2(394) <= r;
scale2(395) <= f_3;
scale2(396) <= f_3;
scale2(397) <= f_3;
scale2(398) <= r;
--------------------25
scale2(399) <= c_3;
scale2(400) <= c_3;
scale2(401) <= c_3;
scale2(402) <= r;
scale2(403) <= am_3;
scale2(404) <= am_3;
scale2(405) <= am_3;
scale2(406) <= am_3;
scale2(407) <= r;
scale2(408) <= r;
scale2(409) <= am_4;
scale2(410) <= am_4;
scale2(411) <= am_4;
scale2(412) <= am_4;
scale2(413) <= r;
scale2(414) <= r;
--------------------26
scale2(415) <= c_4;
scale2(416) <= c_4;
scale2(417) <= c_4;
scale2(418) <= c_4;
scale2(419) <= r;
scale2(420) <= r;
scale2(421) <= g_3;
scale2(422) <= r;
scale2(423) <= g_3;
scale2(424) <= g_3;
scale2(425) <= g_3;
scale2(426) <= r;
scale2(427) <= c_3;
scale2(428) <= c_3;
scale2(429) <= c_3;
scale2(430) <= r;
--------------------27
scale2(431) <= am_2;
scale2(432) <= am_2;
scale2(433) <= am_2;
scale2(434) <= am_2;
scale2(435) <= r;
scale2(436) <= r;
scale2(437) <= em_4;
scale2(438) <= em_4;
scale2(439) <= r;
scale2(440) <= r;
scale2(441) <= r;
scale2(442) <= r;
scale2(443) <= am_3;
scale2(444) <= am_3;
scale2(445) <= am_3;
scale2(446) <= r;
--------------------28
scale2(447) <= g_3;
scale2(448) <= g_3;
scale2(449) <= g_3;
scale2(450) <= g_3;
scale2(451) <= r;
scale2(452) <= r;
scale2(453) <= c_3;
scale2(454) <= c_3;
scale2(455) <= r;
scale2(456) <= r;
scale2(457) <= r;
scale2(458) <= r;
scale2(459) <= g_2;
scale2(460) <= g_2;
scale2(461) <= g_2;
scale2(462) <= g_2;
--------------------29
scale2(463) <= am_2;
scale2(464) <= am_2;
scale2(465) <= am_2;
scale2(466) <= am_2;
scale2(467) <= r;
scale2(468) <= r;
scale2(469) <= em_4;
scale2(470) <= em_4;
scale2(471) <= r;
scale2(472) <= r;
scale2(473) <= r;
scale2(474) <= r;
scale2(475) <= am_3;
scale2(476) <= am_3;
scale2(477) <= am_3;
scale2(478) <= r;
--------------------30
scale2(479) <= g_3;
scale2(480) <= g_3;
scale2(481) <= g_3;
scale2(482) <= g_3;
scale2(483) <= r;
scale2(484) <= r;
scale2(485) <= c_3;
scale2(486) <= c_3;
scale2(487) <= r;
scale2(488) <= r;
scale2(489) <= r;
scale2(490) <= r;
scale2(491) <= g_2;
scale2(492) <= g_2;
scale2(493) <= g_2;
scale2(494) <= g_2;
--------------------31
scale2(495) <= am_2;
scale2(496) <= am_2;
scale2(497) <= am_2;
scale2(498) <= am_2;
scale2(499) <= r;
scale2(500) <= r;
scale2(501) <= em_4;
scale2(502) <= em_4;
scale2(503) <= r;
scale2(504) <= r;
scale2(505) <= r;
scale2(506) <= r;
scale2(507) <= am_3;
scale2(508) <= am_3;
scale2(509) <= am_3;
scale2(510) <= r;
--------------------32
scale2(511) <= g_3;
scale2(512) <= g_3;
scale2(513) <= g_3;
scale2(514) <= g_3;
scale2(515) <= r;
scale2(516) <= r;
scale2(517) <= c_3;
scale2(518) <= c_3;
scale2(519) <= r;
scale2(520) <= r;
scale2(521) <= r;
scale2(522) <= r;
scale2(523) <= g_2;
scale2(524) <= g_2;
scale2(525) <= g_2;
scale2(526) <= g_2;
--------------------33
scale2(527) <= d_3;
scale2(528) <= r;
scale2(529) <= d_3;
scale2(530) <= d_3;
scale2(531) <= r;
scale2(532) <= r;
scale2(533) <= d_3;
scale2(534) <= d_3;
scale2(535) <= r;
scale2(536) <= r;
scale2(537) <= d_3;
scale2(538) <= r;
scale2(539) <= d_3;
scale2(540) <= d_3;
scale2(541) <= d_3;
scale2(542) <= r;
--------------------34
scale2(543) <= g_3;
scale2(544) <= g_3;
scale2(545) <= g_3;
scale2(546) <= g_3;
scale2(547) <= r;
scale2(548) <= r;
scale2(549) <= r;
scale2(550) <= r;
scale2(551) <= g_2;
scale2(552) <= g_2;
scale2(553) <= g_2;
scale2(554) <= g_2;
scale2(555) <= r;
scale2(556) <= r;
scale2(557) <= r;
scale2(558) <= r;
-----2---------------35
scale2(559) <= g_3;
scale2(560) <= g_3;
scale2(561) <= g_3;
scale2(562) <= g_3;
scale2(563) <= r;
scale2(564) <= r;
scale2(565) <= e_3;
scale2(566) <= e_3;
scale2(567) <= e_3;
scale2(568) <= e_3;
scale2(569) <= r;
scale2(570) <= r;
scale2(571) <= c_3;
scale2(572) <= c_3;
scale2(573) <= c_3;
scale2(574) <= c_3;
-----2---------------36
scale2(575) <= r;
scale2(576) <= r;
scale2(577) <= f_3;
scale2(578) <= f_3;
scale2(579) <= f_3;
scale2(580) <= r;
scale2(581) <= g_3;
scale2(582) <= g_3;
scale2(583) <= g_3;
scale2(584) <= r;
scale2(585) <= gm_3;
scale2(586) <= r;
scale2(587) <= f_3;
scale2(588) <= f_3;
scale2(589) <= f_3;
scale2(590) <= r;
-----2---------------37
scale2(591) <= e_3;
scale2(592) <= e_3;
scale2(593) <= r;
scale2(594) <= c_4;
scale2(595) <= c_4;
scale2(596) <= r;
scale2(597) <= e_4;
scale2(598) <= r;
scale2(599) <= f_4;
scale2(600) <= f_4;
scale2(601) <= f_4;
scale2(602) <= r;
scale2(603) <= d_4;
scale2(604) <= r;
scale2(605) <= e_4;
scale2(606) <= e_4;
-----2---------------38
scale2(607) <= r;
scale2(608) <= r;
scale2(609) <= c_4;
scale2(610) <= c_4;
scale2(611) <= c_4;
scale2(612) <= r;
scale2(613) <= a_4;
scale2(614) <= r;
scale2(615) <= b_4;
scale2(616) <= r;
scale2(617) <= g_4;
scale2(618) <= g_4;
scale2(619) <= g_4;
scale2(620) <= g_4;
scale2(621) <= r;
scale2(622) <= r;
-----2---------------39
scale2(623) <= g_3;
scale2(624) <= g_3;
scale2(625) <= g_3;
scale2(626) <= g_3;
scale2(627) <= r;
scale2(628) <= r;
scale2(629) <= e_3;
scale2(630) <= e_3;
scale2(631) <= e_3;
scale2(632) <= e_3;
scale2(633) <= r;
scale2(634) <= r;
scale2(635) <= c_3;
scale2(636) <= c_3;
scale2(637) <= c_3;
scale2(638) <= c_3;
-----2---------------40
scale2(639) <= r;
scale2(640) <= r;
scale2(641) <= f_3;
scale2(642) <= f_3;
scale2(643) <= f_3;
scale2(644) <= r;
scale2(645) <= g_3;
scale2(646) <= g_3;
scale2(647) <= g_3;
scale2(648) <= r;
scale2(649) <= gm_3;
scale2(650) <= r;
scale2(651) <= f_3;
scale2(652) <= f_3;
scale2(653) <= f_3;
scale2(654) <= r;
-----2---------------41
scale2(655) <= e_3;
scale2(656) <= e_3;
scale2(657) <= r;
scale2(658) <= c_4;
scale2(659) <= c_4;
scale2(660) <= r;
scale2(661) <= e_4;
scale2(662) <= r;
scale2(663) <= f_4;
scale2(664) <= f_4;
scale2(665) <= f_4;
scale2(666) <= r;
scale2(667) <= d_4;
scale2(668) <= r;
scale2(669) <= e_4;
scale2(670) <= e_4;
-----2---------------42
scale2(671) <= r;
scale2(672) <= r;
scale2(673) <= c_4;
scale2(674) <= c_4;
scale2(675) <= c_4;
scale2(676) <= r;
scale2(677) <= a_4;
scale2(678) <= r;
scale2(679) <= b_4;
scale2(680) <= r;
scale2(681) <= g_4;
scale2(682) <= g_4;
scale2(683) <= g_4;
scale2(684) <= g_4;
scale2(685) <= r;
scale2(686) <= r;
-----2---------------43
scale2(687) <= c_3;
scale2(688) <= c_3;
scale2(689) <= c_3;
scale2(690) <= c_3;
scale2(691) <= r;
scale2(692) <= r;
scale2(693) <= gm_3;
scale2(694) <= r;
scale2(695) <= g_3;
scale2(696) <= g_3;
scale2(697) <= g_3;
scale2(698) <= r;
scale2(699) <= c_4;
scale2(700) <= c_4;
scale2(701) <= c_4;
scale2(702) <= r;
-----2---------------44
scale2(703) <= f_3;
scale2(704) <= f_3;
scale2(705) <= f_3;
scale2(706) <= r;
scale2(707) <= f_3;
scale2(708) <= f_3;
scale2(709) <= f_3;
scale2(710) <= r;
scale2(711) <= c_4;
scale2(712) <= r;
scale2(713) <= c_4;
scale2(714) <= r;
scale2(715) <= f_3;
scale2(716) <= f_3;
scale2(717) <= f_3;
scale2(718) <= r;
-----2---------------45
scale2(719) <= d_3;
scale2(720) <= d_3;
scale2(721) <= d_3;
scale2(722) <= d_3;
scale2(723) <= r;
scale2(724) <= r;
scale2(725) <= f_3;
scale2(726) <= r;
scale2(727) <= g_3;
scale2(728) <= g_3;
scale2(729) <= g_3;
scale2(730) <= r;
scale2(731) <= b_4;
scale2(732) <= b_4;
scale2(733) <= b_4;
scale2(734) <= r;
-----2---------------46
scale2(735) <= g_3;
scale2(736) <= g_3;
scale2(737) <= g_3;
scale2(738) <= r;
scale2(739) <= g_3;
scale2(740) <= g_3;
scale2(741) <= g_3;
scale2(742) <= r;
scale2(743) <= c_4;
scale2(744) <= r;
scale2(745) <= c_4;
scale2(746) <= r;
scale2(747) <= g_3;
scale2(748) <= g_3;
scale2(749) <= g_3;
scale2(750) <= r;
-----2---------------47
scale2(751) <= c_3;
scale2(752) <= c_3;
scale2(753) <= c_3;
scale2(754) <= c_3;
scale2(755) <= r;
scale2(756) <= r;
scale2(757) <= gm_3;
scale2(758) <= r;
scale2(759) <= g_3;
scale2(760) <= g_3;
scale2(761) <= g_3;
scale2(762) <= r;
scale2(763) <= c_4;
scale2(764) <= c_4;
scale2(765) <= c_4;
scale2(766) <= r;
-----2---------------48
scale2(767) <= f_3;
scale2(768) <= f_3;
scale2(769) <= f_3;
scale2(770) <= r;
scale2(771) <= f_3;
scale2(772) <= f_3;
scale2(773) <= f_3;
scale2(774) <= r;
scale2(775) <= c_4;
scale2(776) <= r;
scale2(777) <= c_4;
scale2(778) <= r;
scale2(779) <= f_3;
scale2(780) <= f_3;
scale2(781) <= f_3;
scale2(782) <= r;
-----2---------------49
scale2(783) <= g_3;
scale2(784) <= r;
scale2(785) <= g_3;
scale2(786) <= g_3;
scale2(787) <= g_3;
scale2(788) <= r;
scale2(789) <= g_3;
scale2(790) <= r;
scale2(791) <= g_3;
scale2(792) <= g_3;
scale2(793) <= r;
scale2(794) <= a_4;
scale2(795) <= a_4;
scale2(796) <= r; 
scale2(797) <= b_4;
scale2(798) <= r;
-----2--------------50
scale2(799) <= c_4;
scale2(800) <= c_4;
scale2(801) <= c_4;
scale2(802) <= r;
scale2(803) <= g_3;
scale2(804) <= g_3;
scale2(805) <= g_3;
scale2(806) <= r;
scale2(807) <= c_3;
scale2(808) <= c_3;
scale2(809) <= c_3;
scale2(810) <= c_3;
scale2(811) <= r;
scale2(812) <= r;
scale2(813) <= r;
scale2(814) <= r;
-----2-------------51
scale2(815) <= c_3;
scale2(816) <= c_3;
scale2(817) <= c_3;
scale2(818) <= c_3;
scale2(819) <= r;
scale2(820) <= r;
scale2(821) <= gm_3;
scale2(822) <= r;
scale2(823) <= g_3;
scale2(824) <= g_3;
scale2(825) <= g_3;
scale2(826) <= r;
scale2(827) <= c_4;
scale2(828) <= c_4;
scale2(829) <= c_4;
scale2(830) <= r;
-----2--------------52
scale2(831) <= f_3;
scale2(832) <= f_3;
scale2(833) <= f_3;
scale2(834) <= r;
scale2(835) <= f_3;
scale2(836) <= f_3;
scale2(837) <= f_3;
scale2(838) <= r;
scale2(839) <= c_4;
scale2(840) <= r;
scale2(841) <= c_4;
scale2(842) <= r;
scale2(843) <= f_3;
scale2(844) <= f_3;
scale2(845) <= f_3;
scale2(846) <= r;
-----2--------------53
scale2(847) <= d_3;
scale2(848) <= d_3;
scale2(849) <= d_3;
scale2(850) <= d_3;
scale2(851) <= r;
scale2(852) <= r;
scale2(853) <= f_3;
scale2(854) <= r;
scale2(855) <= g_3;
scale2(856) <= g_3;
scale2(857) <= g_3;
scale2(858) <= r;
scale2(859) <= b_4;
scale2(860) <= b_4;
scale2(861) <= b_4;
scale2(862) <= r;
--------------------54
scale2(863) <= g_3;
scale2(864) <= g_3;
scale2(865) <= g_3;
scale2(866) <= r;
scale2(867) <= g_3;
scale2(868) <= g_3;
scale2(869) <= g_3;
scale2(870) <= r;
scale2(871) <= c_4;
scale2(872) <= r;
scale2(873) <= c_4;
scale2(874) <= r;
scale2(875) <= g_3;
scale2(876) <= g_3;
scale2(877) <= g_3;
scale2(878) <= r;
-----2---------------55
scale2(879) <= c_3;
scale2(880) <= c_3;
scale2(881) <= c_3;
scale2(882) <= c_3;
scale2(883) <= r;
scale2(884) <= r;
scale2(885) <= gm_3;
scale2(886) <= r;
scale2(887) <= g_3;
scale2(888) <= g_3;
scale2(889) <= g_3;
scale2(890) <= r;
scale2(891) <= c_4;
scale2(892) <= c_4;
scale2(893) <= c_4;
scale2(894) <= r;
-----2---------------56
scale2(895) <= f_3;
scale2(896) <= f_3;
scale2(897) <= f_3;
scale2(898) <= r;
scale2(899) <= f_3;
scale2(900) <= f_3;
scale2(901) <= f_3;
scale2(902) <= r;
scale2(903) <= c_4;
scale2(904) <= r;
scale2(905) <= c_4;
scale2(906) <= r;
scale2(907) <= f_3;
scale2(908) <= f_3;
scale2(909) <= f_3;
scale2(910) <= r;
-----2--------------57
scale2(911) <= g_3;
scale2(912) <= r;
scale2(913) <= g_3;
scale2(914) <= g_3;
scale2(915) <= g_3;
scale2(916) <= r;
scale2(917) <= g_3;
scale2(918) <= r;
scale2(919) <= g_3;
scale2(920) <= g_3;
scale2(921) <= r;
scale2(922) <= a_4;
scale2(923) <= a_4;
scale2(924) <= r; 
scale2(925) <= b_4;
scale2(926) <= r;
-----2--------------58
scale2(927) <= c_4;
scale2(928) <= c_4;
scale2(929) <= c_4;
scale2(930) <= r;
scale2(931) <= g_3;
scale2(932) <= g_3;
scale2(933) <= g_3;
scale2(934) <= r;
scale2(935) <= c_3;
scale2(936) <= c_3;
scale2(937) <= c_3;
scale2(938) <= c_3;
scale2(939) <= r;
scale2(940) <= r;
scale2(941) <= r;
scale2(942) <= r;
-----2--------------59
scale2(943) <= am_2;
scale2(944) <= am_2;
scale2(945) <= am_2;
scale2(946) <= am_2;
scale2(947) <= r;
scale2(948) <= r;
scale2(949) <= em_4;
scale2(950) <= em_4;
scale2(951) <= r;
scale2(952) <= r;
scale2(953) <= r;
scale2(954) <= r;
scale2(955) <= am_3;
scale2(956) <= am_3;
scale2(957) <= am_3;
scale2(958) <= r;
------------------60
scale2(959) <= g_3;
scale2(960) <= g_3;
scale2(961) <= g_3;
scale2(962) <= g_3;
scale2(963) <= r;
scale2(964) <= r;
scale2(965) <= c_3;
scale2(966) <= c_3;
scale2(967) <= r;
scale2(968) <= r;
scale2(969) <= r;
scale2(970) <= r;
scale2(971) <= g_2;
scale2(972) <= g_2;
scale2(973) <= g_2;
scale2(974) <= g_2;
-----2-------------61
scale2(975) <= am_2;
scale2(976) <= am_2;
scale2(977) <= am_2;
scale2(978) <= am_2;
scale2(979) <= r;
scale2(980) <= r;
scale2(981) <= em_4;
scale2(982) <= em_4;
scale2(983) <= r;
scale2(984) <= r;
scale2(985) <= r;
scale2(986) <= r;
scale2(987) <= am_3;
scale2(988) <= am_3;
scale2(989) <= am_3;
scale2(990) <= r;
-----2---------------62
scale2(991) <= g_3;
scale2(992) <= g_3;
scale2(993) <= g_3;
scale2(994) <= g_3;
scale2(995) <= r;
scale2(996) <= r;
scale2(997) <= c_3;
scale2(998) <= c_3;
scale2(999) <= r;
scale2(1000) <= r;
scale2(1001) <= r;
scale2(1002) <= r;
scale2(1003) <= g_2;
scale2(1004) <= g_2;
scale2(1005) <= g_2;
scale2(1006) <= g_2;
-----2---------------63
scale2(1007) <= am_2;
scale2(1008) <= am_2;
scale2(1009) <= am_2;
scale2(1010) <= am_2;
scale2(1011) <= r;
scale2(1012) <= r;
scale2(1013) <= em_4;
scale2(1014) <= em_4;
scale2(1015) <= r;
scale2(1016) <= r;
scale2(1017) <= r;
scale2(1018) <= r;
scale2(1019) <= am_3;
scale2(1020) <= am_3;
scale2(1021) <= am_3;
scale2(1022) <= r;
-----2---------------64
scale2(1023) <= g_3;
scale2(1024) <= g_3;
scale2(1025) <= g_3;
scale2(1026) <= g_3;
scale2(1027) <= r;
scale2(1028) <= r;
scale2(1029) <= c_3;
scale2(1030) <= c_3;
scale2(1031) <= r;
scale2(1032) <= r;
scale2(1033) <= r;
scale2(1034) <= r;
scale2(1035) <= g_2;
scale2(1036) <= g_2;
scale2(1037) <= g_2;
scale2(1038) <= g_2;
-----2---------------65
scale2(1039) <= d_3;
scale2(1040) <= r;
scale2(1041) <= d_3;
scale2(1042) <= d_3;
scale2(1043) <= r;
scale2(1044) <= r;
scale2(1045) <= d_3;
scale2(1046) <= d_3;
scale2(1047) <= r;
scale2(1048) <= r;
scale2(1049) <= d_3;
scale2(1050) <= r;
scale2(1051) <= d_3;
scale2(1052) <= d_3;
scale2(1053) <= d_3;
scale2(1054) <= r;
-----2---------------66
scale2(1055) <= g_3;
scale2(1056) <= g_3;
scale2(1057) <= g_3;
scale2(1058) <= g_3;
scale2(1059) <= r;
scale2(1060) <= r;
scale2(1061) <= r;
scale2(1062) <= r;
scale2(1063) <= g_2;
scale2(1064) <= g_2;
scale2(1065) <= g_2;
scale2(1066) <= g_2;
scale2(1067) <= r;
scale2(1068) <= r;
scale2(1069) <= r;
scale2(1070) <= r;
-----2---------------67
scale2(1071) <= c_3;
scale2(1072) <= c_3;
scale2(1073) <= c_3;
scale2(1074) <= c_3;
scale2(1075) <= r;
scale2(1076) <= r;
scale2(1077) <= gm_3;
scale2(1078) <= r;
scale2(1079) <= g_3;
scale2(1080) <= g_3;
scale2(1081) <= g_3;
scale2(1082) <= r;
scale2(1083) <= c_4;
scale2(1084) <= c_4;
scale2(1085) <= c_4;
scale2(1086) <= r;
--------------------68
scale2(1087) <= f_3;
scale2(1088) <= f_3;
scale2(1089) <= f_3;
scale2(1090) <= r;
scale2(1091) <= f_3;
scale2(1092) <= f_3;
scale2(1093) <= f_3;
scale2(1094) <= r;
scale2(1095) <= c_4;
scale2(1096) <= r;
scale2(1097) <= c_4;
scale2(1098) <= r;
scale2(1099) <= f_3;
scale2(1100) <= f_3;
scale2(1101) <= f_3;
scale2(1102) <= r;
-----2---------------69
scale2(1103) <= d_3;
scale2(1104) <= d_3;
scale2(1105) <= d_3;
scale2(1106) <= d_3;
scale2(1107) <= r;
scale2(1108) <= r;
scale2(1109) <= f_3;
scale2(1110) <= r;
scale2(1111) <= g_3;
scale2(1112) <= g_3;
scale2(1113) <= g_3;
scale2(1114) <= r;
scale2(1115) <= b_4;
scale2(1116) <= b_4;
scale2(1117) <= b_4;
scale2(1118) <= r;
-----2---------------70
scale2(1119) <= g_3;
scale2(1120) <= g_3;
scale2(1121) <= g_3;
scale2(1122) <= r;
scale2(1123) <= g_3;
scale2(1124) <= g_3;
scale2(1125) <= g_3;
scale2(1126) <= r;
scale2(1127) <= c_4;
scale2(1128) <= r;
scale2(1129) <= c_4;
scale2(1130) <= r;
scale2(1131) <= g_3;
scale2(1132) <= g_3;
scale2(1133) <= g_3;
scale2(1134) <= r;
-----2---------------71
scale2(1135) <= c_3;
scale2(1136) <= c_3;
scale2(1137) <= c_3;
scale2(1138) <= c_3;
scale2(1139) <= r;
scale2(1140) <= r;
scale2(1141) <= gm_3;
scale2(1142) <= r;
scale2(1143) <= g_3;
scale2(1144) <= g_3;
scale2(1145) <= g_3;
scale2(1146) <= r;
scale2(1147) <= c_4;
scale2(1148) <= c_4;
scale2(1149) <= c_4;
scale2(1150) <= r;
------22--------------72
scale2(1151) <= f_3;
scale2(1152) <= f_3;
scale2(1153) <= f_3;
scale2(1154) <= r;
scale2(1155) <= f_3;
scale2(1156) <= f_3;
scale2(1157) <= f_3;
scale2(1158) <= r;
scale2(1159) <= c_4;
scale2(1160) <= r;
scale2(1161) <= c_4;
scale2(1162) <= r;
scale2(1163) <= f_3;
scale2(1164) <= f_3;
scale2(1165) <= f_3;
scale2(1166) <= r;
-----2---------------73
scale2(1167) <= g_3;
scale2(1168) <= r;
scale2(1169) <= g_3;
scale2(1170) <= g_3;
scale2(1171) <= g_3;
scale2(1172) <= r;
scale2(1173) <= g_3;
scale2(1174) <= r;
scale2(1175) <= g_3;
scale2(1176) <= g_3;
scale2(1177) <= r;
scale2(1178) <= a_4;
scale2(1179) <= a_4;
scale2(1180) <= r; 
scale2(1181) <= b_4;
scale2(1182) <= r;
-----2---------------74
scale2(1183) <= c_4;
scale2(1184) <= c_4;
scale2(1185) <= c_4;
scale2(1186) <= r;
scale2(1187) <= g_3;
scale2(1188) <= g_3;
scale2(1189) <= g_3;
scale2(1190) <= r;
scale2(1191) <= c_3;
scale2(1192) <= c_3;
scale2(1193) <= c_3;
scale2(1194) <= c_3;
scale2(1195) <= r;
scale2(1196) <= r;
scale2(1197) <= r;
scale2(1198) <= r;
-----2---------------75
scale2(1199) <= c_3;
scale2(1200) <= c_3;
scale2(1201) <= c_3;
scale2(1202) <= c_3;
scale2(1203) <= r;
scale2(1204) <= r;
scale2(1205) <= gm_3;
scale2(1206) <= r;
scale2(1207) <= g_3;
scale2(1208) <= g_3;
scale2(1209) <= g_3;
scale2(1210) <= r;
scale2(1211) <= c_4;
scale2(1212) <= c_4;
scale2(1213) <= c_4;
scale2(1214) <= r;
-----2---------------76
scale2(1215) <= f_3;
scale2(1216) <= f_3;
scale2(1217) <= f_3;
scale2(1218) <= r;
scale2(1219) <= f_3;
scale2(1220) <= f_3;
scale2(1221) <= f_3;
scale2(1222) <= r;
scale2(1223) <= c_4;
scale2(1224) <= r;
scale2(1225) <= c_4;
scale2(1226) <= r;
scale2(1227) <= f_3;
scale2(1228) <= f_3;
scale2(1229) <= f_3;
scale2(1230) <= r;
-----2---------------77
scale2(1231) <= d_3;
scale2(1232) <= d_3;
scale2(1233) <= d_3;
scale2(1234) <= d_3;
scale2(1235) <= r;
scale2(1236) <= r;
scale2(1237) <= f_3;
scale2(1238) <= r;
scale2(1239) <= g_3;
scale2(1240) <= g_3;
scale2(1241) <= g_3;
scale2(1242) <= r;
scale2(1243) <= b_4;
scale2(1244) <= b_4;
scale2(1245) <= b_4;
scale2(1246) <= r;
-----2---------------78
scale2(1247) <= g_3;
scale2(1248) <= g_3;
scale2(1249) <= g_3;
scale2(1250) <= r;
scale2(1251) <= g_3;
scale2(1252) <= g_3;
scale2(1253) <= g_3;
scale2(1254) <= r;
scale2(1255) <= c_4;
scale2(1256) <= r;
scale2(1257) <= c_4;
scale2(1258) <= r;
scale2(1259) <= g_3;
scale2(1260) <= g_3;
scale2(1261) <= g_3;
scale2(1262) <= r;
-----2---------------79
scale2(1263) <= c_3;
scale2(1264) <= c_3;
scale2(1265) <= c_3;
scale2(1266) <= c_3;
scale2(1267) <= r;
scale2(1268) <= r;
scale2(1269) <= gm_3;
scale2(1270) <= r;
scale2(1271) <= g_3;
scale2(1272) <= g_3;
scale2(1273) <= g_3;
scale2(1274) <= r;
scale2(1275) <= c_4;
scale2(1276) <= c_4;
scale2(1277) <= c_4;
scale2(1278) <= r;
-----2---------------80
scale2(1279) <= f_3;
scale2(1280) <= f_3;
scale2(1281) <= f_3;
scale2(1282) <= r;
scale2(1283) <= f_3;
scale2(1284) <= f_3;
scale2(1285) <= f_3;
scale2(1286) <= r;
scale2(1287) <= c_4;
scale2(1288) <= r;
scale2(1289) <= c_4;
scale2(1290) <= r;
scale2(1291) <= f_3;
scale2(1292) <= f_3;
scale2(1293) <= f_3;
scale2(1294) <= r;
-----2---------------81
scale2(1295) <= g_3;
scale2(1296) <= r;
scale2(1297) <= g_3;
scale2(1298) <= g_3;
scale2(1299) <= g_3;
scale2(1300) <= r;
scale2(1301) <= g_3;
scale2(1302) <= r;
scale2(1303) <= g_3;
scale2(1304) <= g_3;
scale2(1305) <= r;
scale2(1306) <= a_4;
scale2(1307) <= a_4;
scale2(1308) <= r; 
scale2(1309) <= b_4;
scale2(1310) <= r;
-----2---------------82
scale2(1311) <= c_4;
scale2(1312) <= c_4;
scale2(1313) <= c_4;
scale2(1314) <= r;
scale2(1315) <= g_3;
scale2(1316) <= g_3;
scale2(1317) <= g_3;
scale2(1318) <= r;
scale2(1319) <= c_3;
scale2(1320) <= c_3;
scale2(1321) <= c_3;
scale2(1322) <= c_3;
scale2(1323) <= r;
scale2(1324) <= r;
scale2(1325) <= r;
scale2(1326) <= r;
-----2---------------83
scale2(1327) <= g_3;
scale2(1328) <= g_3;
scale2(1329) <= g_3;
scale2(1330) <= g_3;
scale2(1331) <= r;
scale2(1332) <= r;
scale2(1333) <= e_3;
scale2(1334) <= e_3;
scale2(1335) <= e_3;
scale2(1336) <= e_3;
scale2(1337) <= r;
scale2(1338) <= r;
scale2(1339) <= c_3;
scale2(1340) <= c_3;
scale2(1341) <= c_3;
scale2(1342) <= r;
-----2---------------84
scale2(1343) <= c_3;
scale2(1344) <= c_3;
scale2(1345) <= c_3;
scale2(1346) <= c_3;
scale2(1347) <= c_3;
scale2(1348) <= c_3;
scale2(1349) <= c_3;
scale2(1350) <= r;
scale2(1351) <= am_2;
scale2(1352) <= am_2;
scale2(1353) <= am_2;
scale2(1354) <= am_2;
scale2(1355) <= am_2;
scale2(1356) <= am_2;
scale2(1357) <= am_2;
scale2(1358) <= r;
-----2---------------85
scale2(1359) <= g_2;
scale2(1360) <= g_2;
scale2(1361) <= g_2;
scale2(1362) <= g_2;
scale2(1363) <= g_2;
scale2(1364) <= g_2;
scale2(1365) <= g_2;
scale2(1366) <= g_2;
scale2(1367) <= g_2;
scale2(1368) <= g_2;
scale2(1369) <= g_2;
scale2(1370) <= g_2;
scale2(1371) <= g_2;
scale2(1372) <= g_2;
scale2(1373) <= g_2;
scale2(1374) <= g_2;


		

process (n_clk,rss,rst)
begin
   if rss = '1' or rst = '1' then
      dot_data_00 <= zr;
		dot_data_01 <= zr;
		dot_data_02 <= zr;
		dot_data_03 <= zr;
		dot_data_04 <= zr;
		dot_data_05 <= zr;
		dot_data_06 <= zr;
		dot_data_07 <= zr;
		dot_data_08 <= zr;
		dot_data_09 <= zr;
		dot_data_10 <= zr;
		dot_data_11 <= zr;
		dot_data_12 <= zr;
		dot_data_13 <= zr;
		d_dp <= zr;
		d_d  <= zr;
		d_dm <= zr;		
	elsif n_clk'event and n_clk = '1' then
		d_dp        <= dot_data_00;
		d_d         <= dot_data_01;
		d_dm        <= dot_data_02;
		dot_data_00 <= dot_data_01;
		dot_data_01 <= dot_data_02;
		dot_data_02 <= dot_data_03;
		dot_data_03 <= dot_data_04;
		dot_data_04 <= dot_data_05;
		dot_data_05 <= dot_data_06;
		dot_data_06 <= dot_data_07;
		dot_data_07 <= dot_data_08;
		dot_data_08 <= dot_data_09;
		dot_data_09 <= dot_data_10;
		dot_data_10 <= dot_data_11;
		dot_data_11 <= dot_data_12;
		dot_data_12 <= dot_data_13;
		dot_data_13 <= data_b(note);
	end if;
end process;




u0 : dot_dis
port map (
	clk => clk,
	dot_data_00 => dot_data_00,
	dot_data_01 => dot_data_01,
	dot_data_02 => dot_data_02,
	dot_data_03 => dot_data_03,
	dot_data_04 => dot_data_04,
	dot_data_05 => dot_data_05,
	dot_data_06 => dot_data_06,
	dot_data_07 => dot_data_07,
	dot_data_08 => dot_data_08,
	dot_data_09 => dot_data_09,
	dot_data_10 => dot_data_10,
	dot_data_11 => dot_data_11,
	dot_data_12 => dot_data_12,
	dot_data_13 => dot_data_13,
	dot_d => dot_d,
	dot_scan => dot_scan 
);
----------------------------------------------------------------piezo
-------------dot + 15
scale(0) <= r;
scale(1) <= r;
scale(2) <= r;
scale(3) <= r;
scale(4) <= r;
scale(5) <= r;
scale(6) <= r;
scale(7) <= r;
scale(8) <= r;
scale(9) <= r;
scale(10) <= r;
scale(11) <= r;
scale(12) <= r;
scale(13) <= r;
scale(14) <= r;
--------------------1
scale(15) <= e_5;
scale(16) <= r;
scale(17) <= e_5;
scale(18) <= e_5;
scale(19) <= r;
scale(20) <= r;
scale(21) <= e_5;
scale(22) <= e_5;
scale(23) <= r;
scale(24) <= r;
scale(25) <= c_5;
scale(26) <= r;
scale(27) <= e_5;
scale(28) <= e_5;
scale(29) <= e_5;
scale(30) <= r;
-------------------2
scale(31) <= g_5;
scale(32) <= g_5;
scale(33) <= g_5;
scale(34) <= g_5;
scale(35) <= r;
scale(36) <= r;
scale(37) <= r;
scale(38) <= r;
scale(39) <= g_4;
scale(40) <= g_4;
scale(41) <= g_4;
scale(42) <= g_4;
scale(43) <= r;
scale(44) <= r;
scale(45) <= r;
scale(46) <= r;
-------------------3
scale(47) <= c_5;
scale(48) <= c_5;
scale(49) <= c_5;
scale(50) <= c_5;
scale(51) <= r;
scale(52) <= r;
scale(53) <= g_4;
scale(54) <= g_4;
scale(55) <= g_4;
scale(56) <= g_4;
scale(57) <= r;
scale(58) <= r;
scale(59) <= e_4;
scale(60) <= e_4;
scale(61) <= e_4;
scale(62) <= e_4;
-------------------4
scale(63) <= r;
scale(64) <= r;
scale(65) <= a_5;
scale(66) <= a_5;
scale(67) <= a_5;
scale(68) <= r;
scale(69) <= b_5;
scale(70) <= b_5;
scale(71) <= b_5;
scale(72) <= r;
scale(73) <= bm_5;
scale(74) <= bm_5;
scale(75) <= a_5;
scale(76) <= a_5;
scale(77) <= a_5;
scale(78) <= r;
--------------------5
scale(79) <= g_4;
scale(80) <= g_4;
scale(81) <= r;
scale(82) <= e_5;
scale(83) <= e_5;
scale(84) <= r;
scale(85) <= g_5;
scale(86) <= r;
scale(87) <= a_6;
scale(88) <= a_6;
scale(89) <= a_6;
scale(90) <= r;
scale(91) <= f_5;
scale(92) <= r;
scale(93) <= g_5;
scale(94) <= g_5;
--------------------6
scale(95) <= r;
scale(96) <= r;
scale(97) <= e_5;
scale(98) <= e_5;
scale(99) <= e_5;
scale(100) <= r;
scale(101) <= c_5;
scale(102) <= r;
scale(103) <= d_5;
scale(104) <= r;
scale(105) <= b_5;
scale(106) <= b_5;
scale(107) <= b_5;
scale(108) <= b_5;
scale(109) <= r;
scale(110) <= r;
--------------------7
scale(111) <= c_5;
scale(112) <= c_5;
scale(113) <= c_5;
scale(114) <= c_5;
scale(115) <= r;
scale(116) <= r;
scale(117) <= g_4;
scale(118) <= g_4;
scale(119) <= g_4;
scale(120) <= g_4;
scale(121) <= r;
scale(122) <= r;
scale(123) <= e_4;
scale(124) <= e_4;
scale(125) <= e_4;
scale(126) <= e_4;
-----------------------8
scale(127) <= r;
scale(128) <= r;
scale(129) <= a_5;
scale(130) <= a_5;
scale(131) <= a_5;
scale(132) <= r;
scale(133) <= b_5;
scale(134) <= b_5;
scale(135) <= b_5;
scale(136) <= r;
scale(137) <= bm_5;
scale(138) <= r;
scale(139) <= a_5;
scale(140) <= a_5;
scale(141) <= a_5;
scale(142) <= r;
----------------------9
scale(143) <= g_4;
scale(144) <= g_4;
scale(145) <= r;
scale(146) <= e_5;
scale(147) <= e_5;
scale(148) <= r;
scale(149) <= g_5;
scale(150) <= r;
scale(151) <= a_6;
scale(152) <= a_6;
scale(153) <= a_6;
scale(154) <= r;
scale(155) <= f_5;
scale(156) <= r;
scale(157) <= g_5;
scale(158) <= g_5;
---------------------10
scale(159) <= r;
scale(160) <= r;
scale(161) <= e_5;
scale(162) <= e_5;
scale(163) <= e_5;
scale(164) <= r;
scale(165) <= c_5;
scale(166) <= r;
scale(167) <= d_5;
scale(168) <= r;
scale(169) <= b_5;
scale(170) <= b_5;
scale(171) <= b_5;
scale(172) <= b_5;
scale(173) <= r;
scale(174) <= r;
---------------------11
scale(175) <= r;
scale(176) <= r;
scale(177) <= r;
scale(178) <= r;
scale(179) <= g_5;
scale(180) <= r;
scale(181) <= gm_5;
scale(182) <= r;
scale(183) <= f_5;
scale(184) <= r;
scale(185) <= em_5;
scale(186) <= em_5;
scale(187) <= em_5;
scale(188) <= r;
scale(189) <= e_5;
scale(190) <= e_5;
---------------------12
scale(191) <= r;
scale(192) <= r;
scale(193) <= am_4;
scale(194) <= r;
scale(195) <= a_5;
scale(196) <= r;
scale(197) <= c_5;
scale(198) <= c_5;
scale(199) <= r;
scale(200) <= r;
scale(201) <= a_5;
scale(202) <= r;
scale(203) <= c_5;
scale(204) <= r;
scale(205) <= d_5;
scale(206) <= d_5;
---------------------13
scale(207) <= r;
scale(208) <= r;
scale(209) <= r;
scale(210) <= r;
scale(211) <= g_5;
scale(212) <= r;
scale(213) <= gm_5;
scale(214) <= r;
scale(215) <= f_5;
scale(216) <= r;
scale(217) <= em_5;
scale(218) <= em_5;
scale(219) <= em_5;
scale(220) <= r;
scale(221) <= e_5;
scale(222) <= e_5;
---------------------14
scale(223) <= r;
scale(224) <= r;
scale(225) <= c_6;
scale(226) <= c_6;
scale(227) <= c_6;
scale(228) <= r;
scale(229) <= c_6;
scale(230) <= r;
scale(231) <= c_6;
scale(232) <= c_6;
scale(233) <= c_6;
scale(234) <= c_6;
scale(235) <= r;
scale(236) <= r;
scale(237) <= r;
scale(238) <= r;
---------------------15
scale(239) <= r;
scale(240) <= r;
scale(241) <= r;
scale(242) <= r;
scale(243) <= g_5;
scale(244) <= r;
scale(245) <= gm_5;
scale(246) <= r;
scale(247) <= f_5;
scale(248) <= r;
scale(249) <= em_5;
scale(250) <= em_5;
scale(251) <= em_5;
scale(252) <= r;
scale(253) <= e_5;
scale(254) <= e_5;
--------------------16
scale(255) <= r;
scale(256) <= r;
scale(257) <= am_4;
scale(258) <= r;
scale(259) <= a_5;
scale(260) <= r;
scale(261) <= c_5;
scale(262) <= c_5;
scale(263) <= r;
scale(264) <= r;
scale(265) <= a_5;
scale(266) <= r;
scale(267) <= c_5;
scale(268) <= r;
scale(269) <= d_5;
scale(270) <= d_5;
---------------------17
scale(271) <= r;
scale(272) <= r;
scale(273) <= r;
scale(274) <= r;
scale(275) <= em_5;
scale(276) <= em_5;
scale(277) <= em_5;
scale(278) <= em_5;
scale(279) <= r;
scale(280) <= r;
scale(281) <= d_5;
scale(282) <= d_5;
scale(283) <= d_5;
scale(284) <= d_5;
scale(285) <= r;
scale(286) <= r;
--------------------18
scale(287) <= c_5;
scale(288) <= c_5;
scale(289) <= c_5;
scale(290) <= c_5;
scale(291) <= r;
scale(292) <= r;
scale(293) <= r;
scale(294) <= r;
scale(295) <= r;
scale(296) <= r;
scale(297) <= r;
scale(298) <= r;
scale(299) <= r;
scale(300) <= r;
scale(301) <= r;
scale(302) <= r;
---------------------19
scale(303) <= r;
scale(304) <= r;
scale(305) <= r;
scale(306) <= r;
scale(307) <= g_5;
scale(308) <= r;
scale(309) <= gm_5;
scale(310) <= r;
scale(311) <= f_5;
scale(312) <= r;
scale(313) <= em_5;
scale(314) <= em_5;
scale(315) <= em_5;
scale(316) <= r;
scale(317) <= e_5;
scale(318) <= e_5;
--------------------20
scale(319) <= r;
scale(320) <= r;
scale(321) <= am_4;
scale(322) <= r;
scale(323) <= a_5;
scale(324) <= r;
scale(325) <= c_5;
scale(326) <= c_5;
scale(327) <= r;
scale(328) <= r;
scale(329) <= a_5;
scale(330) <= r;
scale(331) <= c_5;
scale(332) <= r;
scale(333) <= d_5;
scale(334) <= d_5;
---------------------21
scale(335) <= r;
scale(336) <= r;
scale(337) <= r;
scale(338) <= r;
scale(339) <= g_5;
scale(340) <= r;
scale(341) <= gm_5;
scale(342) <= r;
scale(343) <= f_5;
scale(344) <= r;
scale(345) <= em_5;
scale(346) <= em_5;
scale(347) <= em_5;
scale(348) <= r;
scale(349) <= e_5;
scale(350) <= e_5;
---------------------22
scale(351) <= r;
scale(352) <= r;
scale(353) <= c_6;
scale(354) <= c_6;
scale(355) <= c_6;
scale(356) <= r;
scale(357) <= c_6;
scale(358) <= r;
scale(359) <= c_6;
scale(360) <= c_6;
scale(361) <= c_6;
scale(362) <= c_6;
scale(363) <= r;
scale(364) <= r;
scale(365) <= r;
scale(366) <= r;
-------------------23
scale(367) <= r;
scale(368) <= r;
scale(369) <= r;
scale(370) <= r;
scale(371) <= g_5;
scale(372) <= r;
scale(373) <= gm_5;
scale(374) <= r;
scale(375) <= f_5;
scale(376) <= r;
scale(377) <= em_5;
scale(378) <= em_5;
scale(379) <= em_5;
scale(380) <= r;
scale(381) <= e_5;
scale(382) <= e_5;
--------------------24
scale(383) <= r;
scale(384) <= r;
scale(385) <= am_4;
scale(386) <= r;
scale(387) <= a_5;
scale(388) <= r;
scale(389) <= c_5;
scale(390) <= c_5;
scale(391) <= r;
scale(392) <= r;
scale(393) <= a_5;
scale(394) <= r;
scale(395) <= c_5;
scale(396) <= r;
scale(397) <= d_5;
scale(398) <= d_5;
---------------------25
scale(399) <= r;
scale(400) <= r;
scale(401) <= r;
scale(402) <= r;
scale(403) <= em_5;
scale(404) <= em_5;
scale(405) <= em_5;
scale(406) <= em_5;
scale(407) <= r;
scale(408) <= r;
scale(409) <= d_5;
scale(410) <= d_5;
scale(411) <= d_5;
scale(412) <= d_5;
scale(413) <= r;
scale(414) <= r;
-------------------26
scale(415) <= c_5;
scale(416) <= c_5;
scale(417) <= c_5;
scale(418) <= c_5;
scale(419) <= r;
scale(420) <= r;
scale(421) <= r;
scale(422) <= r;
scale(423) <= r;
scale(424) <= r;
scale(425) <= r;
scale(426) <= r;
scale(427) <= r;
scale(428) <= r;
scale(429) <= r;
scale(430) <= r;
---------------------27
scale(431) <= c_5;
scale(432) <= r;
scale(433) <= c_5;
scale(434) <= c_5;
scale(435) <= r;
scale(436) <= r;
scale(437) <= c_5;
scale(438) <= c_5;
scale(439) <= r;
scale(440) <= r;
scale(441) <= c_5;
scale(442) <= r;
scale(443) <= d_5;
scale(444) <= d_5;
scale(445) <= d_5;
scale(446) <= r;
--------------------28
scale(447) <= e_5;
scale(448) <= r;
scale(449) <= c_5;
scale(450) <= c_5;
scale(451) <= r;
scale(452) <= r;
scale(453) <= a_5;
scale(454) <= r;
scale(455) <= g_4;
scale(456) <= g_4;
scale(457) <= g_4;
scale(458) <= g_4;
scale(459) <= g_4;
scale(460) <= g_4;
scale(461) <= g_4;
scale(462) <= r;
---------------------29
scale(463) <= c_5;
scale(464) <= r;
scale(465) <= c_5;
scale(466) <= c_5;
scale(467) <= r;
scale(468) <= r;
scale(469) <= c_5;
scale(470) <= c_5;
scale(471) <= r;
scale(472) <= r;
scale(473) <= c_5;
scale(474) <= r;
scale(475) <= d_5;
scale(476) <= r;
scale(477) <= e_5;
scale(478) <= e_5;
-------------------30
scale(479) <= r;
scale(480) <= r;
scale(481) <= r;
scale(482) <= r;
scale(483) <= r;
scale(484) <= r;
scale(485) <= r;
scale(486) <= r;
scale(487) <= r;
scale(488) <= r;
scale(489) <= r;
scale(490) <= r;
scale(491) <= r;
scale(492) <= r;
scale(493) <= r;
scale(494) <= r;
--------------------31
scale(495) <= c_5;
scale(496) <= r;
scale(497) <= c_5;
scale(498) <= c_5;
scale(499) <= r;
scale(500) <= r;
scale(501) <= c_5;
scale(502) <= c_5;
scale(503) <= r;
scale(504) <= r;
scale(505) <= c_5;
scale(506) <= r;
scale(507) <= d_5;
scale(508) <= d_5;
scale(509) <= d_5;
scale(510) <= r;
--------------------32
scale(511) <= e_5;
scale(512) <= r;
scale(513) <= c_5;
scale(514) <= c_5;
scale(515) <= r;
scale(516) <= r;
scale(517) <= a_5;
scale(518) <= r;
scale(519) <= g_4;
scale(520) <= g_4;
scale(521) <= g_4;
scale(522) <= g_4;
scale(523) <= g_4;
scale(524) <= g_4;
scale(525) <= g_4;
scale(526) <= r;
--------------------33
scale(527) <= e_5;
scale(528) <= r;
scale(529) <= e_5;
scale(530) <= e_5;
scale(531) <= r;
scale(532) <= r;
scale(533) <= e_5;
scale(534) <= e_5;
scale(535) <= r;
scale(536) <= r;
scale(537) <= c_5;
scale(538) <= r;
scale(539) <= e_5;
scale(540) <= e_5;
scale(541) <= e_5;
scale(542) <= r;
-------------------34
scale(543) <= g_5;
scale(544) <= g_5;
scale(545) <= g_5;
scale(546) <= g_5;
scale(547) <= r;
scale(548) <= r;
scale(549) <= r;
scale(550) <= r;
scale(551) <= g_4;
scale(552) <= g_4;
scale(553) <= g_4;
scale(554) <= g_4;
scale(555) <= r;
scale(556) <= r;
scale(557) <= r;
scale(558) <= r;
-------------------35
scale(559) <= c_5;
scale(560) <= c_5;
scale(561) <= c_5;
scale(562) <= c_5;
scale(563) <= r;
scale(564) <= r;
scale(565) <= g_4;
scale(566) <= g_4;
scale(567) <= g_4;
scale(568) <= g_4;
scale(569) <= r;
scale(570) <= r;
scale(571) <= e_4;
scale(572) <= e_4;
scale(573) <= e_4;
scale(574) <= e_4;
-------------------36
scale(575) <= r;
scale(576) <= r;
scale(577) <= a_5;
scale(578) <= a_5;
scale(579) <= a_5;
scale(580) <= r;
scale(581) <= b_5;
scale(582) <= b_5;
scale(583) <= b_5;
scale(584) <= r;
scale(585) <= bm_5;
scale(586) <= bm_5;
scale(587) <= a_5;
scale(588) <= a_5;
scale(589) <= a_5;
scale(590) <= r;
--------------------37
scale(591) <= g_4;
scale(592) <= g_4;
scale(593) <= r;
scale(594) <= e_5;
scale(595) <= e_5;
scale(596) <= r;
scale(597) <= g_5;
scale(598) <= r;
scale(599) <= a_6;
scale(600) <= a_6;
scale(601) <= a_6;
scale(602) <= r;
scale(603) <= f_5;
scale(604) <= r;
scale(605) <= g_5;
scale(606) <= g_5;
--------------------38
scale(607) <= r;
scale(608) <= r;
scale(609) <= e_5;
scale(610) <= e_5;
scale(611) <= e_5;
scale(612) <= r;
scale(613) <= c_5;
scale(614) <= r;
scale(615) <= d_5;
scale(616) <= r;
scale(617) <= b_5;
scale(618) <= b_5;
scale(619) <= b_5;
scale(620) <= b_5;
scale(621) <= r;
scale(622) <= r;
--------------------39
scale(623) <= c_5;
scale(624) <= c_5;
scale(625) <= c_5;
scale(626) <= c_5;
scale(627) <= r;
scale(628) <= r;
scale(629) <= g_4;
scale(630) <= g_4;
scale(631) <= g_4;
scale(632) <= g_4;
scale(633) <= r;
scale(634) <= r;
scale(635) <= e_4;
scale(636) <= e_4;
scale(637) <= e_4;
scale(638) <= e_4;
----------------------40
scale(639) <= r;
scale(640) <= r;
scale(641) <= a_5;
scale(642) <= a_5;
scale(643) <= a_5;
scale(644) <= r;
scale(645) <= b_5;
scale(646) <= b_5;
scale(647) <= b_5;
scale(648) <= r;
scale(649) <= bm_5;
scale(650) <= r;
scale(651) <= a_5;
scale(652) <= a_5;
scale(653) <= a_5;
scale(654) <= r;
--------------------41
scale(655) <= g_4;
scale(656) <= g_4;
scale(657) <= r;
scale(658) <= e_5;
scale(659) <= e_5;
scale(660) <= r;
scale(661) <= g_5;
scale(662) <= r;
scale(663) <= a_6;
scale(664) <= a_6;
scale(665) <= a_6;
scale(666) <= r;
scale(667) <= f_5;
scale(668) <= r;
scale(669) <= g_5;
scale(670) <= g_5;
-------------------42
scale(671) <= r;
scale(672) <= r;
scale(673) <= e_5;
scale(674) <= e_5;
scale(675) <= e_5;
scale(676) <= r;
scale(677) <= c_5;
scale(678) <= r;
scale(679) <= d_5;
scale(680) <= r;
scale(681) <= b_5;
scale(682) <= b_5;
scale(683) <= b_5;
scale(684) <= b_5;
scale(685) <= r;
scale(686) <= r;
--------------------43
scale(687) <= e_5;
scale(688) <= r;
scale(689) <= c_5;
scale(690) <= c_5;
scale(691) <= c_5;
scale(692) <= r;
scale(693) <= g_4;
scale(694) <= g_4;
scale(695) <= r;
scale(696) <= r;
scale(697) <= r;
scale(698) <= r;
scale(699) <= am_4;
scale(700) <= am_4;
scale(701) <= am_4;
scale(702) <= r;
--------------------44
scale(703) <= a_5;
scale(704) <= r;
scale(705) <= f_5;
scale(706) <= f_5;
scale(707) <= f_5;
scale(708) <= r;
scale(709) <= f_5;
scale(710) <= r;
scale(711) <= a_5;
scale(712) <= a_5;
scale(713) <= a_5;
scale(714) <= a_5;
scale(715) <= r;
scale(716) <= r;
scale(717) <= r;
scale(718) <= r;
-------------------45
scale(719) <= b_5;
scale(720) <= b_5;
scale(721) <= r;
scale(722) <= a_6;
scale(723) <= a_6;
scale(724) <= r;
scale(725) <= a_6;
scale(726) <= r;
scale(727) <= a_6;
scale(728) <= a_6;
scale(729) <= r;
scale(730) <= g_5;
scale(731) <= g_5;
scale(732) <= r;
scale(733) <= f_5;
scale(734) <= r;
------------------46
scale(735) <= e_5;
scale(736) <= r;
scale(737) <= c_5;
scale(738) <= c_5;
scale(739) <= c_5;
scale(740) <= r;
scale(741) <= a_5;
scale(742) <= r;
scale(743) <= g_4;
scale(744) <= g_4;
scale(745) <= g_4;
scale(746) <= g_4;
scale(747) <= r;
scale(748) <= r;
scale(749) <= r;
scale(750) <= r;
--------------------47
scale(751) <= e_5;
scale(752) <= r;
scale(753) <= c_5;
scale(754) <= c_5;
scale(755) <= c_5;
scale(756) <= r;
scale(757) <= g_4;
scale(758) <= g_4;
scale(759) <= r;
scale(760) <= r;
scale(761) <= r;
scale(762) <= r;
scale(763) <= am_4;
scale(764) <= am_4;
scale(765) <= am_4;
scale(766) <= r;
------------------48
scale(767) <= a_5;
scale(768) <= r;
scale(769) <= f_5;
scale(770) <= f_5;
scale(771) <= f_5;
scale(772) <= r;
scale(773) <= f_5;
scale(774) <= r;
scale(775) <= a_5;
scale(776) <= a_5;
scale(777) <= a_5;
scale(778) <= a_5;
scale(779) <= r;
scale(780) <= r;
scale(781) <= r;
scale(782) <= r;
--------------------49
scale(783) <= b_5;
scale(784) <= r;
scale(785) <= f_5;
scale(786) <= f_5;
scale(787) <= f_5;
scale(788) <= r;
scale(789) <= f_5;
scale(790) <= r;
scale(791) <= f_5;
scale(792) <= f_5;
scale(793) <= r;
scale(794) <= e_5;
scale(795) <= e_5;
scale(796) <= r;
scale(797) <= d_5;
scale(798) <= r;
--------------------50
scale(799) <= c_5;
scale(800) <= r;
scale(801) <= e_4;
scale(802) <= e_4;
scale(803) <= e_4;
scale(804) <= r;
scale(805) <= e_4;
scale(806) <= r;
scale(807) <= c_4;
scale(808) <= c_4;
scale(809) <= c_4;
scale(810) <= c_4;
scale(811) <= r;
scale(812) <= r;
scale(813) <= r;
scale(814) <= r;
----------------------51
scale(815) <= e_5;
scale(816) <= r;
scale(817) <= c_5;
scale(818) <= c_5;
scale(819) <= c_5;
scale(820) <= r;
scale(821) <= g_4;
scale(822) <= g_4;
scale(823) <= r;
scale(824) <= r;
scale(825) <= r;
scale(826) <= r;
scale(827) <= am_4;
scale(828) <= am_4;
scale(829) <= am_4;
scale(830) <= r;
-------------------52
scale(831) <= a_5;
scale(832) <= r;
scale(833) <= f_5;
scale(834) <= f_5;
scale(835) <= f_5;
scale(836) <= r;
scale(837) <= f_5;
scale(838) <= r;
scale(839) <= a_5;
scale(840) <= a_5;
scale(841) <= a_5;
scale(842) <= a_5;
scale(843) <= r;
scale(844) <= r;
scale(845) <= r;
scale(846) <= r;
-------------------53
scale(847) <= b_5;
scale(848) <= b_5;
scale(849) <= r;
scale(850) <= a_6;
scale(851) <= a_6;
scale(852) <= r;
scale(853) <= a_6;
scale(854) <= r;
scale(855) <= a_6;
scale(856) <= a_6;
scale(857) <= r;
scale(858) <= g_5;
scale(859) <= g_5;
scale(860) <= r;
scale(861) <= f_5;
scale(862) <= r;
---------------------54
scale(863) <= e_5;
scale(864) <= r;
scale(865) <= c_5;
scale(866) <= c_5;
scale(867) <= c_5;
scale(868) <= r;
scale(869) <= a_5;
scale(870) <= r;
scale(871) <= g_4;
scale(872) <= g_4;
scale(873) <= g_4;
scale(874) <= g_4;
scale(875) <= r;
scale(876) <= r;
scale(877) <= r;
scale(878) <= r;
---------------------55
scale(879) <= e_5;
scale(880) <= r;
scale(881) <= c_5;
scale(882) <= c_5;
scale(883) <= c_5;
scale(884) <= r;
scale(885) <= g_4;
scale(886) <= g_4;
scale(887) <= r;
scale(888) <= r;
scale(889) <= r;
scale(890) <= r;
scale(891) <= am_4;
scale(892) <= am_4;
scale(893) <= am_4;
scale(894) <= r;
------------------56
scale(895) <= a_5;
scale(896) <= r;
scale(897) <= f_5;
scale(898) <= f_5;
scale(899) <= f_5;
scale(900) <= r;
scale(901) <= f_5;
scale(902) <= r;
scale(903) <= a_5;
scale(904) <= a_5;
scale(905) <= a_5;
scale(906) <= a_5;
scale(907) <= r;
scale(908) <= r;
scale(909) <= r;
scale(910) <= r;
---------------------57
scale(911) <= b_5;
scale(912) <= r;
scale(913) <= f_5;
scale(914) <= f_5;
scale(915) <= f_5;
scale(916) <= r;
scale(917) <= f_5;
scale(918) <= r;
scale(919) <= f_5;
scale(920) <= f_5;
scale(921) <= r;
scale(922) <= e_5;
scale(923) <= e_5;
scale(924) <= r;
scale(925) <= d_5;
scale(926) <= r;
------------------58
scale(927) <= c_5;
scale(928) <= r;
scale(929) <= e_4;
scale(930) <= e_4;
scale(931) <= e_4;
scale(932) <= r;
scale(933) <= e_4;
scale(934) <= r;
scale(935) <= c_4;
scale(936) <= c_4;
scale(937) <= c_4;
scale(938) <= c_4;
scale(939) <= r;
scale(940) <= r;
scale(941) <= r;
scale(942) <= r;
------------------59
scale(943) <= c_5;
scale(944) <= r;
scale(945) <= c_5;
scale(946) <= c_5;
scale(947) <= r;
scale(948) <= r;
scale(949) <= c_5;
scale(950) <= c_5;
scale(951) <= r;
scale(952) <= r;
scale(953) <= c_5;
scale(954) <= r;
scale(955) <= d_5;
scale(956) <= d_5;
scale(957) <= d_5;
scale(958) <= r;
--------------------60
scale(959) <= e_5;
scale(960) <= r;
scale(961) <= c_5;
scale(962) <= c_5;
scale(963) <= r;
scale(964) <= r;
scale(965) <= a_5;
scale(966) <= r;
scale(967) <= g_4;
scale(968) <= g_4;
scale(969) <= g_4;
scale(970) <= g_4;
scale(971) <= g_4;
scale(972) <= g_4;
scale(973) <= g_4;
scale(974) <= r;
--------------------61
scale(975) <= c_5;
scale(976) <= r;
scale(977) <= c_5;
scale(978) <= c_5;
scale(979) <= r;
scale(980) <= r;
scale(981) <= c_5;
scale(982) <= c_5;
scale(983) <= r;
scale(984) <= r;
scale(985) <= c_5;
scale(986) <= r;
scale(987) <= d_5;
scale(988) <= r;
scale(989) <= e_5;
scale(990) <= e_5;
------------------------62
scale(991) <= r;
scale(992) <= r;
scale(993) <= r;
scale(994) <= r;
scale(995) <= e_5;
scale(996) <= r;
scale(997) <= g_5;
scale(998) <= r;
scale(999) <= e_6;
scale(1000) <= r;
scale(1001) <= c_6;
scale(1002) <= r;
scale(1003) <= d_6;
scale(1004) <= r;
scale(1005) <= g_6;
scale(1006) <= r;
--------------------63
scale(1007) <= c_5;
scale(1008) <= r;
scale(1009) <= c_5;
scale(1010) <= c_5;
scale(1011) <= r;
scale(1012) <= r;
scale(1013) <= c_5;
scale(1014) <= c_5;
scale(1015) <= r;
scale(1016) <= r;
scale(1017) <= c_5;
scale(1018) <= r;
scale(1019) <= d_5;
scale(1020) <= d_5;
scale(1021) <= d_5;
scale(1022) <= r;
--------------------64
scale(1023) <= e_5;
scale(1024) <= r;
scale(1025) <= c_5;
scale(1026) <= c_5;
scale(1027) <= r;
scale(1028) <= r;
scale(1029) <= a_5;
scale(1030) <= r;
scale(1031) <= g_4;
scale(1032) <= g_4;
scale(1033) <= g_4;
scale(1034) <= g_4;
scale(1035) <= g_4;
scale(1036) <= g_4;
scale(1037) <= g_4;
scale(1038) <= r;
---------------------65
scale(1039) <= e_5;
scale(1040) <= r;
scale(1041) <= e_5;
scale(1042) <= e_5;
scale(1043) <= r;
scale(1044) <= r;
scale(1045) <= e_5;
scale(1046) <= e_5;
scale(1047) <= r;
scale(1048) <= r;
scale(1049) <= c_5;
scale(1050) <= r;
scale(1051) <= e_5;
scale(1052) <= e_5;
scale(1053) <= e_5;
scale(1054) <= r;
-------------------66
scale(1055) <= g_5;
scale(1056) <= g_5;
scale(1057) <= g_5;
scale(1058) <= g_5;
scale(1059) <= r;
scale(1060) <= r;
scale(1061) <= r;
scale(1062) <= r;
scale(1063) <= g_4;
scale(1064) <= g_4;
scale(1065) <= g_4;
scale(1066) <= g_4;
scale(1067) <= r;
scale(1068) <= r;
scale(1069) <= r;
scale(1070) <= r;
------------------67
scale(1071) <= e_5;
scale(1072) <= r;
scale(1073) <= c_5;
scale(1074) <= c_5;
scale(1075) <= c_5;
scale(1076) <= r;
scale(1077) <= g_4;
scale(1078) <= g_4;
scale(1079) <= r;
scale(1080) <= r;
scale(1081) <= r;
scale(1082) <= r;
scale(1083) <= am_4;
scale(1084) <= am_4;
scale(1085) <= am_4;
scale(1086) <= r;
--------------------68
scale(1087) <= a_5;
scale(1088) <= r;
scale(1089) <= f_5;
scale(1090) <= f_5;
scale(1091) <= f_5;
scale(1092) <= r;
scale(1093) <= f_5;
scale(1094) <= r;
scale(1095) <= a_5;
scale(1096) <= a_5;
scale(1097) <= a_5;
scale(1098) <= a_5;
scale(1099) <= r;
scale(1100) <= r;
scale(1101) <= r;
scale(1102) <= r;
--------------------69
scale(1103) <= b_5;
scale(1104) <= b_5;
scale(1105) <= r;
scale(1106) <= a_6;
scale(1107) <= a_6;
scale(1108) <= r;
scale(1109) <= a_6;
scale(1110) <= r;
scale(1111) <= a_6;
scale(1112) <= a_6;
scale(1113) <= r;
scale(1114) <= g_5;
scale(1115) <= g_5;
scale(1116) <= r;
scale(1117) <= f_5;
scale(1118) <= r;
--------------------70
scale(1119) <= e_5;
scale(1120) <= r;
scale(1121) <= c_5;
scale(1122) <= c_5;
scale(1123) <= c_5;
scale(1124) <= r;
scale(1125) <= a_5;
scale(1126) <= r;
scale(1127) <= g_4;
scale(1128) <= g_4;
scale(1129) <= g_4;
scale(1130) <= g_4;
scale(1131) <= r;
scale(1132) <= r;
scale(1133) <= r;
scale(1134) <= r;
--------------------71
scale(1135) <= e_5;
scale(1136) <= r;
scale(1137) <= c_5;
scale(1138) <= c_5;
scale(1139) <= c_5;
scale(1140) <= r;
scale(1141) <= g_4;
scale(1142) <= g_4;
scale(1143) <= r;
scale(1144) <= r;
scale(1145) <= r;
scale(1146) <= r;
scale(1147) <= am_4;
scale(1148) <= am_4;
scale(1149) <= am_4;
scale(1150) <= r;
---------------------72
scale(1151) <= a_5;
scale(1152) <= r;
scale(1153) <= f_5;
scale(1154) <= f_5;
scale(1155) <= f_5;
scale(1156) <= r;
scale(1157) <= f_5;
scale(1158) <= r;
scale(1159) <= a_5;
scale(1160) <= a_5;
scale(1161) <= a_5;
scale(1162) <= a_5;
scale(1163) <= r;
scale(1164) <= r;
scale(1165) <= r;
scale(1166) <= r;
---------------------73
scale(1167) <= b_5;
scale(1168) <= r;
scale(1169) <= f_5;
scale(1170) <= f_5;
scale(1171) <= f_5;
scale(1172) <= r;
scale(1173) <= f_5;
scale(1174) <= r;
scale(1175) <= f_5;
scale(1176) <= f_5;
scale(1177) <= r;
scale(1178) <= e_5;
scale(1179) <= e_5;
scale(1180) <= r;
scale(1181) <= d_5;
scale(1182) <= r;
--------------------74
scale(1183) <= c_5;
scale(1184) <= r;
scale(1185) <= e_4;
scale(1186) <= e_4;
scale(1187) <= e_4;
scale(1188) <= r;
scale(1189) <= e_4;
scale(1190) <= r;
scale(1191) <= c_4;
scale(1192) <= c_4;
scale(1193) <= c_4;
scale(1194) <= c_4;
scale(1195) <= r;
scale(1196) <= r;
scale(1197) <= r;
scale(1198) <= r;
------------------75
scale(1199) <= e_5;
scale(1200) <= r;
scale(1201) <= c_5;
scale(1202) <= c_5;
scale(1203) <= c_5;
scale(1204) <= r;
scale(1205) <= g_4;
scale(1206) <= g_4;
scale(1207) <= r;
scale(1208) <= r;
scale(1209) <= r;
scale(1210) <= r;
scale(1211) <= am_4;
scale(1212) <= am_4;
scale(1213) <= am_4;
scale(1214) <= r;
--------------------76
scale(1215) <= a_5;
scale(1216) <= r;
scale(1217) <= f_5;
scale(1218) <= f_5;
scale(1219) <= f_5;
scale(1220) <= r;
scale(1221) <= f_5;
scale(1222) <= r;
scale(1223) <= a_5;
scale(1224) <= a_5;
scale(1225) <= a_5;
scale(1226) <= a_5;
scale(1227) <= r;
scale(1228) <= r;
scale(1229) <= r;
scale(1230) <= r;
--------------------77
scale(1231) <= b_5;
scale(1232) <= b_5;
scale(1233) <= r;
scale(1234) <= a_6;
scale(1235) <= a_6;
scale(1236) <= r;
scale(1237) <= a_6;
scale(1238) <= r;
scale(1239) <= a_6;
scale(1240) <= a_6;
scale(1241) <= r;
scale(1242) <= g_5;
scale(1243) <= g_5;
scale(1244) <= r;
scale(1245) <= f_5;
scale(1246) <= r;
--------------------78
scale(1247) <= e_5;
scale(1248) <= r;
scale(1249) <= c_5;
scale(1250) <= c_5;
scale(1251) <= c_5;
scale(1252) <= r;
scale(1253) <= a_5;
scale(1254) <= r;
scale(1255) <= g_4;
scale(1256) <= g_4;
scale(1257) <= g_4;
scale(1258) <= g_4;
scale(1259) <= r;
scale(1260) <= r;
scale(1261) <= r;
scale(1262) <= r;
-------------------79
scale(1263) <= e_5;
scale(1264) <= r;
scale(1265) <= c_5;
scale(1266) <= c_5;
scale(1267) <= c_5;
scale(1268) <= r;
scale(1269) <= g_4;
scale(1270) <= g_4;
scale(1271) <= r;
scale(1272) <= r;
scale(1273) <= r;
scale(1274) <= r;
scale(1275) <= am_4;
scale(1276) <= am_4;
scale(1277) <= am_4;
scale(1278) <= r;
--------------------80
scale(1279) <= a_5;
scale(1280) <= r;
scale(1281) <= f_5;
scale(1282) <= f_5;
scale(1283) <= f_5;
scale(1284) <= r;
scale(1285) <= f_5;
scale(1286) <= r;
scale(1287) <= a_5;
scale(1288) <= a_5;
scale(1289) <= a_5;
scale(1290) <= a_5;
scale(1291) <= r;
scale(1292) <= r;
scale(1293) <= r;
scale(1294) <= r;
--------------------81
scale(1295) <= b_5;
scale(1296) <= r;
scale(1297) <= f_5;
scale(1298) <= f_5;
scale(1299) <= f_5;
scale(1300) <= r;
scale(1301) <= f_5;
scale(1302) <= r;
scale(1303) <= f_5;
scale(1304) <= f_5;
scale(1305) <= r;
scale(1306) <= e_5;
scale(1307) <= e_5;
scale(1308) <= r;
scale(1309) <= d_5;
scale(1310) <= r;
--------------------82
scale(1311) <= c_5;
scale(1312) <= r;
scale(1313) <= e_4;
scale(1314) <= e_4;
scale(1315) <= e_4;
scale(1316) <= r;
scale(1317) <= e_4;
scale(1318) <= r;
scale(1319) <= c_4;
scale(1320) <= c_4;
scale(1321) <= c_4;
scale(1322) <= c_4;
scale(1323) <= r;
scale(1324) <= r;
scale(1325) <= r;
scale(1326) <= r;
-------------------83
scale(1327) <= c_5;
scale(1328) <= c_5;
scale(1329) <= c_5;
scale(1330) <= c_5;
scale(1331) <= r;
scale(1332) <= r;
scale(1333) <= g_4;
scale(1334) <= g_4;
scale(1335) <= g_4;
scale(1336) <= g_4;
scale(1337) <= r;
scale(1338) <= r;
scale(1339) <= e_4;
scale(1340) <= e_4;
scale(1341) <= e_4;
scale(1342) <= r;
------------------84
scale(1343) <= a_5;
scale(1344) <= a_5;
scale(1345) <= r;
scale(1346) <= b_5;
scale(1347) <= b_5;
scale(1348) <= r;
scale(1349) <= a_5;
scale(1350) <= r;
scale(1351) <= am_4;
scale(1352) <= am_4;
scale(1353) <= r;
scale(1354) <= bm_5;
scale(1355) <= bm_5;
scale(1356) <= r;
scale(1357) <= am_4;
scale(1358) <= r;
-------------------85
scale(1359) <= g_4;
scale(1360) <= g_4;
scale(1361) <= g_4;
scale(1362) <= g_4;
scale(1363) <= g_4;
scale(1364) <= g_4;
scale(1365) <= g_4;
scale(1366) <= g_4;
scale(1367) <= g_4;
scale(1368) <= g_4;
scale(1369) <= g_4;
scale(1370) <= g_4;
scale(1371) <= g_4;
scale(1372) <= g_4;
scale(1373) <= g_4;
scale(1374) <= g_4;
----------------------end

led <= st;

piezo <= p_clk;
piezo2<= p_clk2;
--------------------------------------------------piezo1
process(clk,rst,rss)
begin
  if rst = '1' or rss = '1' then
	  cnt <= 0;
  elsif clk'event and clk = '1' and st = '1' then
     if cnt >= scale(note) then
	     cnt <= 0;
	  else
	     cnt <= cnt + 1;
	  end if;
  end if;
end process;


process (clk,rss,rst)
begin
if rss = '1' or rst = '1' then
  p_clk <= '0';
elsif clk'event and clk = '1' then
	if cnt = 1 then
		p_clk <= not p_clk;
	end if;
end if;
end process;
------------------------------------------------piezo2
process(clk,rst,rss)
begin
  if rst = '1' or rss = '1' then
	  cnt2 <= 0;
  elsif clk'event and clk = '1' and st = '1' then
     if cnt2 >= scale2(note) then
	     cnt2 <= 0;
	  else
	     cnt2 <= cnt2 + 1;
	  end if;
  end if;
end process;


process (clk,rss,rst)
begin
if rss = '1' or rst = '1' then
  p_clk2 <= '0';
elsif clk'event and clk = '1' then
	if cnt2 = 1 then
		p_clk2 <= not p_clk2;
	end if;
end if;
end process;


end a;