----------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

entity mario_hard is
port (
	clk		: in std_logic;     -- 25MHz
	p1       : in std_logic;
	rss      : in std_logic;
	note_clk : out std_logic;
	d_d      : out std_logic_vector(9 downto 0);
	d_dp     : out std_logic_vector(9 downto 0);
	d_dm     : out std_logic_vector(9 downto 0);		
	reset    : out std_logic;	
	rr       : in std_logic;
   -------------------------------------------------------dot port
	dot_d : out std_logic_vector ( 9 downto 0);
	dot_scan : out std_logic_vector ( 13 downto 0);
	--------------------------------------------------------piezo port
	led : out std_logic
);
end mario_hard;

architecture a of mario_hard is
-------------------------------------------------------------------------------component
component dot_dis
port (
	clk : in std_logic;
	dot_data_00 : in std_logic_vector (9 downto 0);
	dot_data_01 : in std_logic_vector (9 downto 0);
	dot_data_02 : in std_logic_vector (9 downto 0);
	dot_data_03 : in std_logic_vector (9 downto 0);
	dot_data_04 : in std_logic_vector (9 downto 0);
	dot_data_05 : in std_logic_vector (9 downto 0);
	dot_data_06 : in std_logic_vector (9 downto 0);
	dot_data_07 : in std_logic_vector (9 downto 0);
	dot_data_08 : in std_logic_vector (9 downto 0);
	dot_data_09 : in std_logic_vector (9 downto 0);
	dot_data_10 : in std_logic_vector (9 downto 0);
	dot_data_11 : in std_logic_vector (9 downto 0);
	dot_data_12 : in std_logic_vector (9 downto 0);
	dot_data_13 : in std_logic_vector (9 downto 0);

	dot_d : out std_logic_vector (9 downto 0);
	dot_scan : out std_logic_vector ( 13 downto 0)
);
end component;
------------------------------------------------------------------------com signal
signal ryt  : integer range 0 to 920312;
signal note : integer range 0 to 1500 := 1450;
signal n_clk   : std_logic := '0';
signal rst : std_logic := '0';

---------------------------------------------------------------------dot signal
signal dot_data_00 : std_logic_vector (9 downto 0);
signal dot_data_01 : std_logic_vector (9 downto 0);
signal dot_data_02 : std_logic_vector (9 downto 0);
signal dot_data_03 : std_logic_vector (9 downto 0);
signal dot_data_04 : std_logic_vector (9 downto 0);
signal dot_data_05 : std_logic_vector (9 downto 0);
signal dot_data_06 : std_logic_vector (9 downto 0);
signal dot_data_07 : std_logic_vector (9 downto 0);
signal dot_data_08 : std_logic_vector (9 downto 0);
signal dot_data_09 : std_logic_vector (9 downto 0);
signal dot_data_10 : std_logic_vector (9 downto 0);
signal dot_data_11 : std_logic_vector (9 downto 0);
signal dot_data_12 : std_logic_vector (9 downto 0);
signal dot_data_13 : std_logic_vector (9 downto 0);

constant zr : std_logic_vector(9 downto 0) := "0000000000";

type data_a is array(1500 downto 0) of std_logic_vector(9 downto 0);
signal data_b : data_a;

--------------------------------------------------------------------piezo signal

signal cnt 	: integer range 0 to 1000000;
signal cnt2 : integer range 0 to 1000000;
signal seq  : integer range 0 to 100000;


signal st   : std_logic := '0';

------------------------------------------------------------------------com

begin

process(p1,rss,rst)
begin
  if p1 = '1' then
     st <= '1';
  elsif rst = '1' or rss = '1' then
     st <= '0';
	  seq <= 0;
  end if;
end process;

process(clk,rst,rss)
begin
  if rst = '1' or rss = '1' then
     ryt <= 0;
	  n_clk <= '0';
  elsif clk'event and clk = '1' and st = '1' then
     if ryt = 920312 then
	     ryt <= 0;
        n_clk <= not n_clk;
     else
        ryt <= ryt + 1;
        n_clk <= n_clk;		  
     end if;
  end if;
end process;

note_clk <= n_clk;

process(n_clk,rss,rst,clk)
begin
  if rss = '1' or rst = '1' then
     note <= 1450;
  elsif n_clk'event and n_clk = '1' then
     if note = 1440 then
	     note <= 1450;
		  rst <= '1';
	  elsif note = 1500 then
	     note <= 0;
	  else
		  note <= note + 1;
     end if;
  end if;
  if rss = '1' or rr = '1' then
     rst <= '0';
  end if;  
end process;

reset <= rst;



---------------------------------------------------------------------dot
data_b(0) <= "0100000001";
data_b(1) <= "0000000000";
data_b(2) <= "0100000001";
data_b(3) <= "0000000000";
data_b(4) <= "0000000000";
data_b(5) <= "0000000000";
data_b(6) <= "0100000001";
data_b(7) <= "0000000000";
data_b(8) <= "0000000000";
data_b(9) <= "0000000000";
data_b(10) <= "0100000010";
data_b(11) <= "0000000000";
data_b(12) <= "0100000001";
data_b(13) <= "0100000001";
data_b(14) <= "0000000000";
data_b(15) <= "0000000000";
--------------------------------1
data_b(16) <= "0001110001";
data_b(17) <= "0001110001";
data_b(18) <= "0000000000";
data_b(19) <= "0000000000";
data_b(20) <= "0000000000";
data_b(21) <= "0000000000";
data_b(22) <= "0000000000";
data_b(23) <= "0000000000";
data_b(24) <= "1000001000";
data_b(25) <= "1000001000";
data_b(26) <= "0000000000";
data_b(27) <= "0000000000";
data_b(28) <= "0000000000";
data_b(29) <= "0000000000";
data_b(30) <= "0000000000";
data_b(31) <= "0000000000";
-----------------------------------2
data_b(32) <= "0001000010";
data_b(33) <= "0001000010";
data_b(34) <= "0000000000";
data_b(35) <= "0000000000";
data_b(36) <= "0000000000";
data_b(37) <= "0000000000";
data_b(38) <= "0010000100";
data_b(39) <= "0010000100";
data_b(40) <= "0000000000";
data_b(41) <= "0000000000";
data_b(42) <= "0000000000";
data_b(43) <= "0000000000";
data_b(44) <= "1000001000";
data_b(45) <= "1000001000";
data_b(46) <= "0000000000";
data_b(47) <= "0000000000";
----------------------------------3
data_b(48) <= "0000000000";
data_b(49) <= "0000000000";
data_b(50) <= "0010001000";
data_b(51) <= "0010001000";
data_b(52) <= "0000000000";
data_b(53) <= "0000000000";
data_b(54) <= "0001000100";
data_b(55) <= "0001000100";
data_b(56) <= "0000000000";
data_b(57) <= "0000000000";
data_b(58) <= "0001000100";
data_b(59) <= "0000000000";
data_b(60) <= "0010001000";
data_b(61) <= "0010001000";
data_b(62) <= "0000000000";
data_b(63) <= "0000000000";
-----------------------------------4
data_b(64) <= "1000001000";
data_b(65) <= "1000001000";
data_b(66) <= "0000000000";
data_b(67) <= "0100000100";
data_b(68) <= "0100000100";
data_b(69) <= "0000000000";
data_b(70) <= "0010000010";
data_b(71) <= "0000000000";
data_b(72) <= "0001000001";
data_b(73) <= "0001000001";
data_b(74) <= "0000000000";
data_b(75) <= "0000000000";
data_b(76) <= "0010000010";
data_b(77) <= "0000000000";
data_b(78) <= "0001000001";
data_b(79) <= "0000000000";
-----------------------------------5
data_b(80) <= "0000000000";
data_b(81) <= "0000000000";
data_b(82) <= "0001000001";
data_b(83) <= "0001000001";
data_b(84) <= "0000000000";
data_b(85) <= "0000000000";
data_b(86) <= "0100000100";
data_b(87) <= "0000000000";
data_b(88) <= "0010000010";
data_b(89) <= "0000000000";
data_b(90) <= "1000001000";
data_b(91) <= "1000001000";
data_b(92) <= "0000000000";
data_b(93) <= "0000000000";
data_b(94) <= "0000000000";
data_b(95) <= "0000000000";
------------------------------------6
data_b(96) <= "0001000010";
data_b(97) <= "0001000010";
data_b(98) <= "0000000000";
data_b(99) <= "0000000000";
data_b(100) <= "0000000000";
data_b(101) <= "0000000000";
data_b(102) <= "0010000100";
data_b(103) <= "0010000100";
data_b(104) <= "0000000000";
data_b(105) <= "0000000000";
data_b(106) <= "0000000000";
data_b(107) <= "0000000000";
data_b(108) <= "1000001000";
data_b(109) <= "1000001000";
data_b(110) <= "0000000000";
data_b(111) <= "0000000000";
----------------------------------7
data_b(112) <= "0000000000";
data_b(113) <= "0000000000";
data_b(114) <= "0010001000";
data_b(115) <= "0010001000";
data_b(116) <= "0000000000";
data_b(117) <= "0000000000";
data_b(118) <= "0001000100";
data_b(119) <= "0001000100";
data_b(120) <= "0000000000";
data_b(121) <= "0000000000";
data_b(122) <= "0001000100";
data_b(123) <= "0000000000";
data_b(124) <= "0010001000";
data_b(125) <= "0010001000";
data_b(126) <= "0000000000";
data_b(127) <= "0000000000";
-----------------------------------8
data_b(128) <= "1000001000";
data_b(129) <= "1000001000";
data_b(130) <= "0000000000";
data_b(131) <= "0100000100";
data_b(132) <= "0100000100";
data_b(133) <= "0000000000";
data_b(134) <= "0010000010";
data_b(135) <= "0000000000";
data_b(136) <= "0001000001";
data_b(137) <= "0001000001";
data_b(138) <= "0000000000";
data_b(139) <= "0000000000";
data_b(140) <= "0010000010";
data_b(141) <= "0000000000";
data_b(142) <= "0001000001";
data_b(143) <= "0000000000";
-----------------------------------9
data_b(144) <= "0000000000";
data_b(145) <= "0000000000";
data_b(146) <= "0001000001";
data_b(147) <= "0001000001";
data_b(148) <= "0000000000";
data_b(149) <= "0000000000";
data_b(150) <= "0100000100";
data_b(151) <= "0000000000";
data_b(152) <= "0010000010";
data_b(153) <= "0000000000";
data_b(154) <= "1000001000";
data_b(155) <= "1000001000";
data_b(156) <= "0000000000";
data_b(157) <= "0000000000";
data_b(158) <= "0000000000";
data_b(159) <= "0000000000";
------------------------------------10
data_b(160) <= "1000000000";
data_b(161) <= "1000000000";
data_b(162) <= "0000000000";
data_b(163) <= "0000000000";
data_b(164) <= "0000000001";
data_b(165) <= "0000000000";
data_b(166) <= "0100000010";
data_b(167) <= "0000000000";
data_b(168) <= "0000000010";
data_b(169) <= "0000000000";
data_b(170) <= "0000001000";
data_b(171) <= "0000001000";
data_b(172) <= "0000000000";
data_b(173) <= "0000000000";
data_b(174) <= "0001000010";
data_b(175) <= "0000000000";
--------------------------------11
data_b(176) <= "0100000000";
data_b(177) <= "0100000000";
data_b(178) <= "0000001000";
data_b(179) <= "0000000000";
data_b(180) <= "0000000100";
data_b(181) <= "0000000000";
data_b(182) <= "0001000010";
data_b(183) <= "0000000000";
data_b(184) <= "0001000000";
data_b(185) <= "0001000000";
data_b(186) <= "0000000100";
data_b(187) <= "0000000000";
data_b(188) <= "0100000010";
data_b(189) <= "0000000000";
data_b(190) <= "0000000001";
data_b(191) <= "0000000000";
----------------------------------12
data_b(192) <= "1000000000";
data_b(193) <= "1000000000";
data_b(194) <= "0000000000";
data_b(195) <= "0000000000";
data_b(196) <= "0000000001";
data_b(197) <= "0000000000";
data_b(198) <= "0100000010";
data_b(199) <= "0000000000";
data_b(200) <= "0000000010";
data_b(201) <= "0000000000";
data_b(202) <= "0000000100";
data_b(203) <= "0000000100";
data_b(204) <= "0010000000";
data_b(205) <= "0000000000";
data_b(206) <= "0001000010";
data_b(207) <= "0000000000";
--------------------------------13
data_b(208) <= "0000000000";
data_b(209) <= "0000000000";
data_b(210) <= "0000110000";
data_b(211) <= "0000110000";
data_b(212) <= "0000000000";
data_b(213) <= "0000000000";
data_b(214) <= "0000110000";
data_b(215) <= "0000000000";
data_b(216) <= "0000110000";
data_b(217) <= "0000110000";
data_b(218) <= "0000000000";
data_b(219) <= "0000000000";
data_b(220) <= "0001000000";
data_b(221) <= "0001000000";
data_b(222) <= "0000000000";
data_b(223) <= "0000000000";
-------------------------------14
data_b(224) <= "1000000000";
data_b(225) <= "1000000000";
data_b(226) <= "0000000000";
data_b(227) <= "0000000000";
data_b(228) <= "0000000001";
data_b(229) <= "0000000000";
data_b(230) <= "0010000010";
data_b(231) <= "0000000000";
data_b(232) <= "0000000010";
data_b(233) <= "0000000000";
data_b(234) <= "0000000100";
data_b(235) <= "0000000100";
data_b(236) <= "0001000000";
data_b(237) <= "0000000000";
data_b(238) <= "0001000010";
data_b(239) <= "0000000000";
-------------------------------15
data_b(240) <= "0100000000";
data_b(241) <= "0100000000";
data_b(242) <= "0100001000";
data_b(243) <= "0000000000";
data_b(244) <= "0000000100";
data_b(245) <= "0000000000";
data_b(246) <= "0001000010";
data_b(247) <= "0000000000";
data_b(248) <= "0001000000";
data_b(249) <= "0001000000";
data_b(250) <= "0001000100";
data_b(251) <= "0000000000";
data_b(252) <= "0100000010";
data_b(253) <= "0100000000";
data_b(254) <= "0100000001";
data_b(255) <= "0100000000";
-----------------------------16
data_b(256) <= "1000000000";
data_b(257) <= "1000000000";
data_b(258) <= "0000000000";
data_b(259) <= "0000000000";
data_b(260) <= "0010000010";
data_b(261) <= "0010000010";
data_b(262) <= "0000000000";
data_b(263) <= "0000000000";
data_b(264) <= "0000000000";
data_b(265) <= "0000000000";
data_b(266) <= "0001000100";
data_b(267) <= "0001000100";
data_b(268) <= "0000000000";
data_b(269) <= "0000000000";
data_b(270) <= "0000000000";
data_b(271) <= "0000000000";
-------------------------------17
data_b(272) <= "0001000100";
data_b(273) <= "0001000100";
data_b(274) <= "0000000000";
data_b(275) <= "0000000000";
data_b(276) <= "0000000000";
data_b(277) <= "0000000000";
data_b(278) <= "0010000000";
data_b(279) <= "0000000000";
data_b(280) <= "0010000000";
data_b(281) <= "0010000000";
data_b(282) <= "0000000000";
data_b(283) <= "0000000000";
data_b(284) <= "1000000000";
data_b(285) <= "1000000000";
data_b(286) <= "0000000000";
data_b(287) <= "0000000000";
--------------------------------18
data_b(288) <= "1000000000";
data_b(289) <= "1000000000";
data_b(290) <= "0000000000";
data_b(291) <= "0000000000";
data_b(292) <= "0000000001";
data_b(293) <= "0000000000";
data_b(294) <= "0100000010";
data_b(295) <= "0000000000";
data_b(296) <= "0000000010";
data_b(297) <= "0000000000";
data_b(298) <= "0000001000";
data_b(299) <= "0000001000";
data_b(300) <= "0000000000";
data_b(301) <= "0000000000";
data_b(302) <= "0001000010";
data_b(303) <= "0000000000";
-------------------------------19
data_b(304) <= "0100000000";
data_b(305) <= "0100000000";
data_b(306) <= "0000001000";
data_b(307) <= "0000000000";
data_b(308) <= "0000000100";
data_b(309) <= "0000000000";
data_b(310) <= "0001000010";
data_b(311) <= "0000000000";
data_b(312) <= "0001000000";
data_b(313) <= "0001000000";
data_b(314) <= "0000000100";
data_b(315) <= "0000000000";
data_b(316) <= "0100000010";
data_b(317) <= "0000000000";
data_b(318) <= "0000000001";
data_b(319) <= "0000000000";
----------------------------------20
data_b(320) <= "1000000000";
data_b(321) <= "1000000000";
data_b(322) <= "0000000000";
data_b(323) <= "0000000000";
data_b(324) <= "0000000001";
data_b(325) <= "0000000000";
data_b(326) <= "0100000010";
data_b(327) <= "0000000000";
data_b(328) <= "0000000010";
data_b(329) <= "0000000000";
data_b(330) <= "0000000100";
data_b(331) <= "0000000100";
data_b(332) <= "0010000000";
data_b(333) <= "0000000000";
data_b(334) <= "0001000010";
data_b(335) <= "0000000000";
--------------------------------21
data_b(336) <= "0000000000";
data_b(337) <= "0000000000";
data_b(338) <= "0000110000";
data_b(339) <= "0000110000";
data_b(340) <= "0000000000";
data_b(341) <= "0000000000";
data_b(342) <= "0000110000";
data_b(343) <= "0000000000";
data_b(344) <= "0000110000";
data_b(345) <= "0000110000";
data_b(346) <= "0000000000";
data_b(347) <= "0000000000";
data_b(348) <= "0001000000";
data_b(349) <= "0001000000";
data_b(350) <= "0000000000";
data_b(351) <= "0000000000";
---------------------------------22
data_b(352) <= "1000000000";
data_b(353) <= "1000000000";
data_b(354) <= "0000000000";
data_b(355) <= "0000000000";
data_b(356) <= "0000000001";
data_b(357) <= "0000000000";
data_b(358) <= "0010000010";
data_b(359) <= "0000000000";
data_b(360) <= "0000000010";
data_b(361) <= "0000000000";
data_b(362) <= "0000000100";
data_b(363) <= "0000000100";
data_b(364) <= "0001000000";
data_b(365) <= "0000000000";
data_b(366) <= "0001000010";
data_b(367) <= "0000000000";
------------------------------23
data_b(368) <= "0100000000";
data_b(369) <= "0100000000";
data_b(370) <= "0100001000";
data_b(371) <= "0000000000";
data_b(372) <= "0000000100";
data_b(373) <= "0000000000";
data_b(374) <= "0001000010";
data_b(375) <= "0000000000";
data_b(376) <= "0001000000";
data_b(377) <= "0001000000";
data_b(378) <= "0001000100";
data_b(379) <= "0000000000";
data_b(380) <= "0100000010";
data_b(381) <= "0100000000";
data_b(382) <= "0100000001";
data_b(383) <= "0100000000";
----------------------------24
data_b(384) <= "1000000000";
data_b(385) <= "1000000000";
data_b(386) <= "0000000000";
data_b(387) <= "0000000000";
data_b(388) <= "0010000010";
data_b(389) <= "0010000010";
data_b(390) <= "0000000000";
data_b(391) <= "0000000000";
data_b(392) <= "0000000000";
data_b(393) <= "0000000000";
data_b(394) <= "0001000100";
data_b(395) <= "0001000100";
data_b(396) <= "0000000000";
data_b(397) <= "0000000000";
data_b(398) <= "0000000000";
data_b(399) <= "0000000000";
----------------------------------25
data_b(400) <= "0001000100";
data_b(401) <= "0001000100";
data_b(402) <= "0000000000";
data_b(403) <= "0000000000";
data_b(404) <= "0000000000";
data_b(405) <= "0000000000";
data_b(406) <= "0010000000";
data_b(407) <= "0000000000";
data_b(408) <= "0010000000";
data_b(409) <= "0010000000";
data_b(410) <= "0000000000";
data_b(411) <= "0000000000";
data_b(412) <= "1000000000";
data_b(413) <= "1000000000";
data_b(414) <= "0000000000";
data_b(415) <= "0000000000";
---------------------------------26
data_b(416) <= "1000000100";
data_b(417) <= "1000000000";
data_b(418) <= "0000000100";
data_b(419) <= "0000000000";
data_b(420) <= "0000000000";
data_b(421) <= "0000000000";
data_b(422) <= "0010000100";
data_b(423) <= "0000000000";
data_b(424) <= "0000000000";
data_b(425) <= "0000000000";
data_b(426) <= "0000000100";
data_b(427) <= "0000000000";
data_b(428) <= "0001000010";
data_b(429) <= "0001000010";
data_b(430) <= "0000000000";
data_b(431) <= "0000000000";
---------------------------------27
data_b(432) <= "0001000001";
data_b(433) <= "0001000000";
data_b(434) <= "0000000010";
data_b(435) <= "0000000000";
data_b(436) <= "0000000000";
data_b(437) <= "0000000000";
data_b(438) <= "0010000100";
data_b(439) <= "0000000000";
data_b(440) <= "0000001000";
data_b(441) <= "0000001000";
data_b(442) <= "0000001000";
data_b(443) <= "0000001000";
data_b(444) <= "1000000000";
data_b(445) <= "1000000000";
data_b(446) <= "0000000000";
data_b(447) <= "0000000000";
------------------------------28
data_b(448) <= "1000000100";
data_b(449) <= "1000000000";
data_b(450) <= "0000000100";
data_b(451) <= "0000000000";
data_b(452) <= "0000000000";
data_b(453) <= "0000000000";
data_b(454) <= "0010000100";
data_b(455) <= "0000000000";
data_b(456) <= "0000000000";
data_b(457) <= "0000000000";
data_b(458) <= "0000000100";
data_b(459) <= "0000000000";
data_b(460) <= "0001000010";
data_b(461) <= "0001000000";
data_b(462) <= "0000000001";
data_b(463) <= "0000000000";
------------------------------29
data_b(464) <= "0001000000";
data_b(465) <= "0001000000";
data_b(466) <= "0000000000";
data_b(467) <= "0000000000";
data_b(468) <= "0000000000";
data_b(469) <= "0000000000";
data_b(470) <= "0010000000";
data_b(471) <= "0000000000";
data_b(472) <= "0000000000";
data_b(473) <= "0000000000";
data_b(474) <= "0000000000";
data_b(475) <= "0000000000";
data_b(476) <= "1000000000";
data_b(477) <= "1000000000";
data_b(478) <= "0000000000";
data_b(479) <= "0000000000";
--------------------------------30
data_b(480) <= "1000000100";
data_b(481) <= "1000000000";
data_b(482) <= "0000000100";
data_b(483) <= "0000000000";
data_b(484) <= "0000000000";
data_b(485) <= "0000000000";
data_b(486) <= "0010000100";
data_b(487) <= "0000000000";
data_b(488) <= "0000000000";
data_b(489) <= "0000000000";
data_b(490) <= "0000000100";
data_b(491) <= "0000000000";
data_b(492) <= "0001000010";
data_b(493) <= "0001000010";
data_b(494) <= "0000000000";
data_b(495) <= "0000000000";
----------------------------------31
data_b(496) <= "0001000001";
data_b(497) <= "0001000000";
data_b(498) <= "0000000010";
data_b(499) <= "0000000000";
data_b(500) <= "0000000000";
data_b(501) <= "0000000000";
data_b(502) <= "0100000100";
data_b(503) <= "0000000000";
data_b(504) <= "0000001000";
data_b(505) <= "0000001000";
data_b(506) <= "0000001000";
data_b(507) <= "0000001000";
data_b(508) <= "1000000000";
data_b(509) <= "1000000000";
data_b(510) <= "0000000000";
data_b(511) <= "0000000000";
----------------------------------32
data_b(512) <= "0100000010";
data_b(513) <= "0000000000";
data_b(514) <= "0100000010";
data_b(515) <= "0000000000";
data_b(516) <= "0000000000";
data_b(517) <= "0000000000";
data_b(518) <= "0100000010";
data_b(519) <= "0000000000";
data_b(520) <= "0000000000";
data_b(521) <= "0000000000";
data_b(522) <= "0100000100";
data_b(523) <= "0000000000";
data_b(524) <= "0100000010";
data_b(525) <= "0100000010";
data_b(526) <= "0000000000";
data_b(527) <= "0000000000";
-----------------------------------33
data_b(528) <= "0001110001";
data_b(529) <= "0001110001";
data_b(530) <= "0000000000";
data_b(531) <= "0000000000";
data_b(532) <= "0000000000";
data_b(533) <= "0000000000";
data_b(534) <= "0000000000";
data_b(535) <= "0000000000";
data_b(536) <= "1000001000";
data_b(537) <= "1000001000";
data_b(538) <= "0000000000";
data_b(539) <= "0000000000";
data_b(540) <= "0000000000";
data_b(541) <= "0000000000";
data_b(542) <= "0000000000";
data_b(543) <= "0000000000";
---------------------------------34
data_b(544) <= "0001000010";
data_b(545) <= "0001000010";
data_b(546) <= "0000000000";
data_b(547) <= "0000000000";
data_b(548) <= "0000000000";
data_b(549) <= "0000000000";
data_b(550) <= "0010000100";
data_b(551) <= "0010000100";
data_b(552) <= "0000000000";
data_b(553) <= "0000000000";
data_b(554) <= "0000000000";
data_b(555) <= "0000000000";
data_b(556) <= "1000001000";
data_b(557) <= "1000001000";
data_b(558) <= "0000000000";
data_b(559) <= "0000000000";
----------------------------------35
data_b(560) <= "0000000000";
data_b(561) <= "0000000000";
data_b(562) <= "0010001000";
data_b(563) <= "0010001000";
data_b(564) <= "0000000000";
data_b(565) <= "0000000000";
data_b(566) <= "0001000100";
data_b(567) <= "0001000100";
data_b(568) <= "0000000000";
data_b(569) <= "0000000000";
data_b(570) <= "0001000100";
data_b(571) <= "0000000000";
data_b(572) <= "0010001000";
data_b(573) <= "0010001000";
data_b(574) <= "0000000000";
data_b(575) <= "0000000000";
----------------------------------36
data_b(576) <= "1000001000";
data_b(577) <= "1000001000";
data_b(578) <= "0000000000";
data_b(579) <= "0100000100";
data_b(580) <= "0100000100";
data_b(581) <= "0000000000";
data_b(582) <= "0010000010";
data_b(583) <= "0000000000";
data_b(584) <= "0001000001";
data_b(585) <= "0001000001";
data_b(586) <= "0000000000";
data_b(587) <= "0000000000";
data_b(588) <= "0010000010";
data_b(589) <= "0000000000";
data_b(590) <= "0001000001";
data_b(591) <= "0000000000";
-----------------------------------37
data_b(592) <= "0000000000";
data_b(593) <= "0000000000";
data_b(594) <= "0001000001";
data_b(595) <= "0001000001";
data_b(596) <= "0000000000";
data_b(597) <= "0000000000";
data_b(598) <= "0100000100";
data_b(599) <= "0000000000";
data_b(600) <= "0010000010";
data_b(601) <= "0000000000";
data_b(602) <= "1000001000";
data_b(603) <= "1000001000";
data_b(604) <= "0000000000";
data_b(605) <= "0000000000";
data_b(606) <= "0000000000";
data_b(607) <= "0000000000";
-----------------------------------38
data_b(608) <= "0001000010";
data_b(609) <= "0001000010";
data_b(610) <= "0000000000";
data_b(611) <= "0000000000";
data_b(612) <= "0000000000";
data_b(613) <= "0000000000";
data_b(614) <= "0010000100";
data_b(615) <= "0010000100";
data_b(616) <= "0000000000";
data_b(617) <= "0000000000";
data_b(618) <= "0000000000";
data_b(619) <= "0000000000";
data_b(620) <= "1000001000";
data_b(621) <= "1000001000";
data_b(622) <= "0000000000";
data_b(623) <= "0000000000";
----------------------------------39
data_b(624) <= "0000000000";
data_b(625) <= "0000000000";
data_b(626) <= "0010001000";
data_b(627) <= "0010001000";
data_b(628) <= "0000000000";
data_b(629) <= "0000000000";
data_b(630) <= "0001000100";
data_b(631) <= "0001000100";
data_b(632) <= "0000000000";
data_b(633) <= "0000000000";
data_b(634) <= "0001000100";
data_b(635) <= "0000000000";
data_b(636) <= "0010001000";
data_b(637) <= "0010001000";
data_b(638) <= "0000000000";
data_b(639) <= "0000000000";
-----------------------------------40
data_b(640) <= "1000001000";
data_b(641) <= "1000001000";
data_b(642) <= "0000000000";
data_b(643) <= "0100000100";
data_b(644) <= "0100000100";
data_b(645) <= "0000000000";
data_b(646) <= "0010000010";
data_b(647) <= "0000000000";
data_b(648) <= "0001000001";
data_b(649) <= "0001000001";
data_b(650) <= "0000000000";
data_b(651) <= "0000000000";
data_b(652) <= "0010000010";
data_b(653) <= "0000000000";
data_b(654) <= "0001000001";
data_b(655) <= "0000000000";
---------------------------------41
data_b(656) <= "0000000000";
data_b(657) <= "0000000000";
data_b(658) <= "0001000001";
data_b(659) <= "0001000001";
data_b(660) <= "0000000000";
data_b(661) <= "0000000000";
data_b(662) <= "0100000100";
data_b(663) <= "0000000000";
data_b(664) <= "0010000010";
data_b(665) <= "0000000000";
data_b(666) <= "1000001000";
data_b(667) <= "1000001000";
data_b(668) <= "0000000000";
data_b(669) <= "0000000000";
data_b(670) <= "0000000000";
data_b(671) <= "0000000000";
-----------------------------------42
data_b(672) <= "1000000001";
data_b(673) <= "1000000000";
data_b(674) <= "0000000010";
data_b(675) <= "0000000000";
data_b(676) <= "0000000000";
data_b(677) <= "0000000000";
data_b(678) <= "0100001000";
data_b(679) <= "0000000000";
data_b(680) <= "0010000000";
data_b(681) <= "0010000000";
data_b(682) <= "0000000000";
data_b(683) <= "0000000000";
data_b(684) <= "0001001000";
data_b(685) <= "0001001000";
data_b(686) <= "0000000000";
data_b(687) <= "0000000000";
------------------------------------43
data_b(688) <= "0100001000";
data_b(689) <= "0100000000";
data_b(690) <= "0000000001";
data_b(691) <= "0000000001";
data_b(692) <= "0100000000";
data_b(693) <= "0100000000";
data_b(694) <= "0000000001";
data_b(695) <= "0000000000";
data_b(696) <= "0001001000";
data_b(697) <= "0000001000";
data_b(698) <= "0001000000";
data_b(699) <= "0000000000";
data_b(700) <= "0100000000";
data_b(701) <= "0100000000";
data_b(702) <= "0000000000";
data_b(703) <= "0000000000";
--------------------------------44
data_b(704) <= "1000001000";
data_b(705) <= "1000001000";
data_b(706) <= "0000000000";
data_b(707) <= "0000000001";
data_b(708) <= "0000000001";
data_b(709) <= "0000000000";
data_b(710) <= "0000000001";
data_b(711) <= "0100000000";
data_b(712) <= "0010000001";
data_b(713) <= "0010000001";
data_b(714) <= "0000000000";
data_b(715) <= "0000000010";
data_b(716) <= "0001000010";
data_b(717) <= "0000000000";
data_b(718) <= "0000000100";
data_b(719) <= "0000000000";
-------------------------------45
data_b(720) <= "0010000001";
data_b(721) <= "0010000000";
data_b(722) <= "0000000010";
data_b(723) <= "0000000010";
data_b(724) <= "0010000000";
data_b(725) <= "0010000000";
data_b(726) <= "0000000100";
data_b(727) <= "0000000000";
data_b(728) <= "0001001000";
data_b(729) <= "0000001000";
data_b(730) <= "0001000000";
data_b(731) <= "0000000000";
data_b(732) <= "0001000000";
data_b(733) <= "0001000000";
data_b(734) <= "0000000000";
data_b(735) <= "0000000000";
-------------------------------46
data_b(736) <= "1000000001";
data_b(737) <= "1000000000";
data_b(738) <= "0000000010";
data_b(739) <= "0000000010";
data_b(740) <= "0000000000";
data_b(741) <= "0000000000";
data_b(742) <= "0100001000";
data_b(743) <= "0000000000";
data_b(744) <= "0010000000";
data_b(745) <= "0010000000";
data_b(746) <= "0000000000";
data_b(747) <= "0000000000";
data_b(748) <= "0001001000";
data_b(749) <= "0001001000";
data_b(750) <= "0000000000";
data_b(751) <= "0000000000";
----------------------------47
data_b(752) <= "0010001000";
data_b(753) <= "0010000000";
data_b(754) <= "0000000001";
data_b(755) <= "0000000001";
data_b(756) <= "0010000000";
data_b(757) <= "0000000000";
data_b(758) <= "0000000001";
data_b(759) <= "0000000000";
data_b(760) <= "0001001000";
data_b(761) <= "0000001000";
data_b(762) <= "0001000000";
data_b(763) <= "0000000000";
data_b(764) <= "0010000000";
data_b(765) <= "0010000000";
data_b(766) <= "0000000000";
data_b(767) <= "0000000000";
--------------------------------48
data_b(768) <= "0100001000";
data_b(769) <= "0000000000";
data_b(770) <= "0100000001";
data_b(771) <= "0100000001";
data_b(772) <= "0000000000";
data_b(773) <= "0000000000";
data_b(774) <= "0100000001";
data_b(775) <= "0000000000";
data_b(776) <= "0100000001";
data_b(777) <= "0100000001";
data_b(778) <= "0000000000";
data_b(779) <= "0010000010";
data_b(780) <= "0010000010";
data_b(781) <= "0000000000";
data_b(782) <= "0001000100";
data_b(783) <= "0000000000";
-------------------------------49
data_b(784) <= "0001000100";
data_b(785) <= "0001000100";
data_b(786) <= "0000000000";
data_b(787) <= "0000000000";
data_b(788) <= "0010000000";
data_b(789) <= "0010000000";
data_b(790) <= "0000000000";
data_b(791) <= "0000000000";
data_b(792) <= "1000000000";
data_b(793) <= "1000000000";
data_b(794) <= "0000000000";
data_b(795) <= "0000000000";
data_b(796) <= "0000000000";
data_b(797) <= "0000000000";
data_b(798) <= "0000000000";
data_b(799) <= "0000000000";
----------------------------50
data_b(800) <= "1000000001";
data_b(801) <= "1000000000";
data_b(802) <= "0000000010";
data_b(803) <= "0000000000";
data_b(804) <= "0000000000";
data_b(805) <= "0000000000";
data_b(806) <= "0100001000";
data_b(807) <= "0000000000";
data_b(808) <= "0010000000";
data_b(809) <= "0010000000";
data_b(810) <= "0000000000";
data_b(811) <= "0000000000";
data_b(812) <= "0001001000";
data_b(813) <= "0001001000";
data_b(814) <= "0000000000";
data_b(815) <= "0000000000";
----------------------------------51
data_b(816) <= "0100001000";
data_b(817) <= "0100000000";
data_b(818) <= "0000000001";
data_b(819) <= "0000000001";
data_b(820) <= "0100000000";
data_b(821) <= "0100000000";
data_b(822) <= "0000000001";
data_b(823) <= "0000000000";
data_b(824) <= "0001001000";
data_b(825) <= "0000001000";
data_b(826) <= "0001000000";
data_b(827) <= "0000000000";
data_b(828) <= "0100000000";
data_b(829) <= "0100000000";
data_b(830) <= "0000000000";
data_b(831) <= "0000000000";
--------------------------------52
data_b(832) <= "1000001000";
data_b(833) <= "1000001000";
data_b(834) <= "0000000000";
data_b(835) <= "0000000001";
data_b(836) <= "0000000001";
data_b(837) <= "0000000000";
data_b(838) <= "0000000001";
data_b(839) <= "0100000000";
data_b(840) <= "0010000001";
data_b(841) <= "0010000001";
data_b(842) <= "0000000000";
data_b(843) <= "0000000010";
data_b(844) <= "0001000010";
data_b(845) <= "0000000000";
data_b(846) <= "0000000100";
data_b(847) <= "0000000000";
------------------------------53
data_b(848) <= "0010000001";
data_b(849) <= "0010000000";
data_b(850) <= "0000000010";
data_b(851) <= "0000000010";
data_b(852) <= "0010000000";
data_b(853) <= "0010000000";
data_b(854) <= "0000000100";
data_b(855) <= "0000000000";
data_b(856) <= "0001001000";
data_b(857) <= "0000001000";
data_b(858) <= "0001000000";
data_b(859) <= "0000000000";
data_b(860) <= "0001000000";
data_b(861) <= "0001000000";
data_b(862) <= "0000000000";
data_b(863) <= "0000000000";
------------------------------54
data_b(864) <= "1000000001";
data_b(865) <= "1000000000";
data_b(866) <= "0000000010";
data_b(867) <= "0000000010";
data_b(868) <= "0000000000";
data_b(869) <= "0000000000";
data_b(870) <= "0100001000";
data_b(871) <= "0000000000";
data_b(872) <= "0010000000";
data_b(873) <= "0010000000";
data_b(874) <= "0000000000";
data_b(875) <= "0000000000";
data_b(876) <= "0001001000";
data_b(877) <= "0001001000";
data_b(878) <= "0000000000";
data_b(879) <= "0000000000";
-----------------------------55
data_b(880) <= "0010001000";
data_b(881) <= "0010000000";
data_b(882) <= "0000000001";
data_b(883) <= "0000000001";
data_b(884) <= "0010000000";
data_b(885) <= "0000000000";
data_b(886) <= "0000000001";
data_b(887) <= "0000000000";
data_b(888) <= "0001001000";
data_b(889) <= "0000001000";
data_b(890) <= "0001000000";
data_b(891) <= "0000000000";
data_b(892) <= "0010000000";
data_b(893) <= "0010000000";
data_b(894) <= "0000000000";
data_b(895) <= "0000000000";
--------------------------------56
data_b(896) <= "0100001000";
data_b(897) <= "0000000000";
data_b(898) <= "0100000001";
data_b(899) <= "0100000001";
data_b(900) <= "0000000000";
data_b(901) <= "0000000000";
data_b(902) <= "0100000001";
data_b(903) <= "0000000000";
data_b(904) <= "0100000001";
data_b(905) <= "0100000001";
data_b(906) <= "0000000000";
data_b(907) <= "0010000010";
data_b(908) <= "0010000010";
data_b(909) <= "0000000000";
data_b(910) <= "0001000100";
data_b(911) <= "0000000000";
-------------------------------57
data_b(912) <= "0001000100";
data_b(913) <= "0001000100";
data_b(914) <= "0000000000";
data_b(915) <= "0000000000";
data_b(916) <= "0010000000";
data_b(917) <= "0010000000";
data_b(918) <= "0000000000";
data_b(919) <= "0000000000";
data_b(920) <= "1000000000";
data_b(921) <= "1000000000";
data_b(922) <= "0000000000";
data_b(923) <= "0000000000";
data_b(924) <= "0000000000";
data_b(925) <= "0000000000";
data_b(926) <= "0000000000";
data_b(927) <= "0000000000";
-----------------------------58
data_b(928) <= "1000000100";
data_b(929) <= "1000000000";
data_b(930) <= "0000000100";
data_b(931) <= "0000000000";
data_b(932) <= "0000000000";
data_b(933) <= "0000000000";
data_b(934) <= "0010000100";
data_b(935) <= "0000000000";
data_b(936) <= "0000000000";
data_b(937) <= "0000000000";
data_b(938) <= "0000000100";
data_b(939) <= "0000000000";
data_b(940) <= "0001000010";
data_b(941) <= "0001000010";
data_b(942) <= "0000000000";
data_b(943) <= "0000000000";
-------------------------------59
data_b(944) <= "0001000001";
data_b(945) <= "0001000000";
data_b(946) <= "0000000010";
data_b(947) <= "0000000000";
data_b(948) <= "0000000000";
data_b(949) <= "0000000000";
data_b(950) <= "0010000100";
data_b(951) <= "0000000000";
data_b(952) <= "0000001000";
data_b(953) <= "0000001000";
data_b(954) <= "0000001000";
data_b(955) <= "0000001000";
data_b(956) <= "1000000000";
data_b(957) <= "1000000000";
data_b(958) <= "0000000000";
data_b(959) <= "0000000000";
-----------------------------60
data_b(960) <= "1000000100";
data_b(961) <= "1000000000";
data_b(962) <= "0000000100";
data_b(963) <= "0000000000";
data_b(964) <= "0000000000";
data_b(965) <= "0000000000";
data_b(966) <= "0010000100";
data_b(967) <= "0000000000";
data_b(968) <= "0000000000";
data_b(969) <= "0000000000";
data_b(970) <= "0000000100";
data_b(971) <= "0000000000";
data_b(972) <= "0001000010";
data_b(973) <= "0001000000";
data_b(974) <= "0000000001";
data_b(975) <= "0000000000";
-------------------------------61
data_b(976) <= "0001000000";
data_b(977) <= "0001000000";
data_b(978) <= "0000000000";
data_b(979) <= "0000000000";
data_b(980) <= "0000001000";
data_b(981) <= "0000000000";
data_b(982) <= "0010000100";
data_b(983) <= "0000000000";
data_b(984) <= "0000110000";
data_b(985) <= "0000000000";
data_b(986) <= "0000000100";
data_b(987) <= "0000000000";
data_b(988) <= "1000000010";
data_b(989) <= "1000000000";
data_b(990) <= "0000110000";
data_b(991) <= "0000000000";
----------------------------62
data_b(992) <= "1000000100";
data_b(993) <= "1000000000";
data_b(994) <= "0000000100";
data_b(995) <= "0000000000";
data_b(996) <= "0000000000";
data_b(997) <= "0000000000";
data_b(998) <= "0010000100";
data_b(999) <= "0000000000";
data_b(1000) <= "0000000000";
data_b(1001) <= "0000000000";
data_b(1002) <= "0000000100";
data_b(1003) <= "0000000000";
data_b(1004) <= "0001000010";
data_b(1005) <= "0001000010";
data_b(1006) <= "0000000000";
data_b(1007) <= "0000000000";
---------------------------------63
data_b(1008) <= "0001000001";
data_b(1009) <= "0001000000";
data_b(1010) <= "0000000010";
data_b(1011) <= "0000000000";
data_b(1012) <= "0000000000";
data_b(1013) <= "0000000000";
data_b(1014) <= "0010000100";
data_b(1015) <= "0000000000";
data_b(1016) <= "0000001000";
data_b(1017) <= "0000001000";
data_b(1018) <= "0000001000";
data_b(1019) <= "0000001000";
data_b(1020) <= "1000000000";
data_b(1021) <= "1000000000";
data_b(1022) <= "0000000000";
data_b(1023) <= "0000000000";
-----------------------------64
data_b(1024) <= "0100000001";
data_b(1025) <= "0000000000";
data_b(1026) <= "0100000001";
data_b(1027) <= "0000000000";
data_b(1028) <= "0000000000";
data_b(1029) <= "0000000000";
data_b(1030) <= "0100000001";
data_b(1031) <= "0000000000";
data_b(1032) <= "0000000000";
data_b(1033) <= "0000000000";
data_b(1034) <= "0100000010";
data_b(1035) <= "0000000000";
data_b(1036) <= "0100000001";
data_b(1037) <= "0100000001";
data_b(1038) <= "0000000000";
data_b(1039) <= "0000000000";
--------------------------------65
data_b(1040) <= "0001110001";
data_b(1041) <= "0001110001";
data_b(1042) <= "0000000000";
data_b(1043) <= "0000000000";
data_b(1044) <= "0000000000";
data_b(1045) <= "0000000000";
data_b(1046) <= "0000000000";
data_b(1047) <= "0000000000";
data_b(1048) <= "1000001000";
data_b(1049) <= "1000001000";
data_b(1050) <= "0000000000";
data_b(1051) <= "0000000000";
data_b(1052) <= "0000000000";
data_b(1053) <= "0000000000";
data_b(1054) <= "0000000000";
data_b(1055) <= "0000000000";
--------------------------------66
data_b(1056) <= "1000000001";
data_b(1057) <= "1000000000";
data_b(1058) <= "0000000010";
data_b(1059) <= "0000000000";
data_b(1060) <= "0000000000";
data_b(1061) <= "0000000000";
data_b(1062) <= "0100001000";
data_b(1063) <= "0000000000";
data_b(1064) <= "0010000000";
data_b(1065) <= "0010000000";
data_b(1066) <= "0000000000";
data_b(1067) <= "0000000000";
data_b(1068) <= "0001001000";
data_b(1069) <= "0001001000";
data_b(1070) <= "0000000000";
data_b(1071) <= "0000000000";
------------------------------------67
data_b(1072) <= "0100001000";
data_b(1073) <= "0100000000";
data_b(1074) <= "0000000001";
data_b(1075) <= "0000000001";
data_b(1076) <= "0100000000";
data_b(1077) <= "0100000000";
data_b(1078) <= "0000000001";
data_b(1079) <= "0000000000";
data_b(1080) <= "0001001000";
data_b(1081) <= "0000001000";
data_b(1082) <= "0001000000";
data_b(1083) <= "0000000000";
data_b(1084) <= "0100000000";
data_b(1085) <= "0100000000";
data_b(1086) <= "0000000000";
data_b(1087) <= "0000000000";
----------------------------------68
data_b(1088) <= "1000001000";
data_b(1089) <= "1000001000";
data_b(1090) <= "0000000000";
data_b(1091) <= "0000000001";
data_b(1092) <= "0000000001";
data_b(1093) <= "0000000000";
data_b(1094) <= "0000000001";
data_b(1095) <= "0100000000";
data_b(1096) <= "0010000001";
data_b(1097) <= "0010000001";
data_b(1098) <= "0000000000";
data_b(1099) <= "0000000010";
data_b(1100) <= "0001000010";
data_b(1101) <= "0000000000";
data_b(1102) <= "0000000100";
data_b(1103) <= "0000000000";
------------------------------69
data_b(1104) <= "0010000001";
data_b(1105) <= "0010000000";
data_b(1106) <= "0000000010";
data_b(1107) <= "0000000010";
data_b(1108) <= "0010000000";
data_b(1109) <= "0010000000";
data_b(1110) <= "0000000100";
data_b(1111) <= "0000000000";
data_b(1112) <= "0001001000";
data_b(1113) <= "0000001000";
data_b(1114) <= "0001000000";
data_b(1115) <= "0000000000";
data_b(1116) <= "0001000000";
data_b(1117) <= "0001000000";
data_b(1118) <= "0000000000";
data_b(1119) <= "0000000000";
--------------------------------70
data_b(1120) <= "1000000001";
data_b(1121) <= "1000000000";
data_b(1122) <= "0000000010";
data_b(1123) <= "0000000010";
data_b(1124) <= "0000000000";
data_b(1125) <= "0000000000";
data_b(1126) <= "0100001000";
data_b(1127) <= "0000000000";
data_b(1128) <= "0010000000";
data_b(1129) <= "0010000000";
data_b(1130) <= "0000000000";
data_b(1131) <= "0000000000";
data_b(1132) <= "0001001000";
data_b(1133) <= "0001001000";
data_b(1134) <= "0000000000";
data_b(1135) <= "0000000000";
-----------------------------71
data_b(1136) <= "0010001000";
data_b(1137) <= "0010000000";
data_b(1138) <= "0000000001";
data_b(1139) <= "0000000001";
data_b(1140) <= "0010000000";
data_b(1141) <= "0000000000";
data_b(1142) <= "0000000001";
data_b(1143) <= "0000000000";
data_b(1144) <= "0001001000";
data_b(1145) <= "0000001000";
data_b(1146) <= "0001000000";
data_b(1147) <= "0000000000";
data_b(1148) <= "0010000000";
data_b(1149) <= "0010000000";
data_b(1150) <= "0000000000";
data_b(1151) <= "0000000000";
---------------------------------72
data_b(1152) <= "0100001000";
data_b(1153) <= "0000000000";
data_b(1154) <= "0100000001";
data_b(1155) <= "0100000001";
data_b(1156) <= "0000000000";
data_b(1157) <= "0000000000";
data_b(1158) <= "0100000001";
data_b(1159) <= "0000000000";
data_b(1160) <= "0100000001";
data_b(1161) <= "0100000001";
data_b(1162) <= "0000000000";
data_b(1163) <= "0010000010";
data_b(1164) <= "0010000010";
data_b(1165) <= "0000000000";
data_b(1166) <= "0001000100";
data_b(1167) <= "0000000000";
--------------------------------73
data_b(1168) <= "0001000100";
data_b(1169) <= "0001000100";
data_b(1170) <= "0000000000";
data_b(1171) <= "0000000000";
data_b(1172) <= "0010000000";
data_b(1173) <= "0010000000";
data_b(1174) <= "0000000000";
data_b(1175) <= "0000000000";
data_b(1176) <= "1000000000";
data_b(1177) <= "1000000000";
data_b(1178) <= "0000000000";
data_b(1179) <= "0000000000";
data_b(1180) <= "0000000000";
data_b(1181) <= "0000000000";
data_b(1182) <= "0000000000";
data_b(1183) <= "0000000000";
-------------------------------------74
data_b(1184) <= "1000000001";
data_b(1185) <= "1000000000";
data_b(1186) <= "0000000010";
data_b(1187) <= "0000000000";
data_b(1188) <= "0000000000";
data_b(1189) <= "0000000000";
data_b(1190) <= "0100001000";
data_b(1191) <= "0000000000";
data_b(1192) <= "0010000000";
data_b(1193) <= "0010000000";
data_b(1194) <= "0000000000";
data_b(1195) <= "0000000000";
data_b(1196) <= "0001001000";
data_b(1197) <= "0001001000";
data_b(1198) <= "0000000000";
data_b(1199) <= "0000000000";
-------------------------------------75
data_b(1200) <= "0100001000";
data_b(1201) <= "0100000000";
data_b(1202) <= "0000000001";
data_b(1203) <= "0000000001";
data_b(1204) <= "0100000000";
data_b(1205) <= "0100000000";
data_b(1206) <= "0000000001";
data_b(1207) <= "0000000000";
data_b(1208) <= "0001001000";
data_b(1209) <= "0000001000";
data_b(1210) <= "0001000000";
data_b(1211) <= "0000000000";
data_b(1212) <= "0100000000";
data_b(1213) <= "0100000000";
data_b(1214) <= "0000000000";
data_b(1215) <= "0000000000";
----------------------------------76
data_b(1216) <= "1000001000";
data_b(1217) <= "1000001000";
data_b(1218) <= "0000000000";
data_b(1219) <= "0000000001";
data_b(1220) <= "0000000001";
data_b(1221) <= "0000000000";
data_b(1222) <= "0000000001";
data_b(1223) <= "0100000000";
data_b(1224) <= "0010000001";
data_b(1225) <= "0010000001";
data_b(1226) <= "0000000000";
data_b(1227) <= "0000000010";
data_b(1228) <= "0001000010";
data_b(1229) <= "0000000000";
data_b(1230) <= "0000000100";
data_b(1231) <= "0000000000";
-------------------------------77
data_b(1232) <= "0010000001";
data_b(1233) <= "0010000000";
data_b(1234) <= "0000000010";
data_b(1235) <= "0000000010";
data_b(1236) <= "0010000000";
data_b(1237) <= "0010000000";
data_b(1238) <= "0000000100";
data_b(1239) <= "0000000000";
data_b(1240) <= "0001001000";
data_b(1241) <= "0000001000";
data_b(1242) <= "0001000000";
data_b(1243) <= "0000000000";
data_b(1244) <= "0001000000";
data_b(1245) <= "0001000000";
data_b(1246) <= "0000000000";
data_b(1247) <= "0000000000";
-------------------------------78
data_b(1248) <= "1000000001";
data_b(1249) <= "1000000000";
data_b(1250) <= "0000000010";
data_b(1251) <= "0000000010";
data_b(1252) <= "0000000000";
data_b(1253) <= "0000000000";
data_b(1254) <= "0100001000";
data_b(1255) <= "0000000000";
data_b(1256) <= "0010000000";
data_b(1257) <= "0010000000";
data_b(1258) <= "0000000000";
data_b(1259) <= "0000000000";
data_b(1260) <= "0001001000";
data_b(1261) <= "0001001000";
data_b(1262) <= "0000000000";
data_b(1263) <= "0000000000";
-----------------------------79
data_b(1264) <= "0010001000";
data_b(1265) <= "0010000000";
data_b(1266) <= "0000000001";
data_b(1267) <= "0000000001";
data_b(1268) <= "0010000000";
data_b(1269) <= "0000000000";
data_b(1270) <= "0000000001";
data_b(1271) <= "0000000000";
data_b(1272) <= "0001001000";
data_b(1273) <= "0000001000";
data_b(1274) <= "0001000000";
data_b(1275) <= "0000000000";
data_b(1276) <= "0010000000";
data_b(1277) <= "0010000000";
data_b(1278) <= "0000000000";
data_b(1279) <= "0000000000";
----------------------------------80
data_b(1280) <= "0100001000";
data_b(1281) <= "0000000000";
data_b(1282) <= "0100000001";
data_b(1283) <= "0100000001";
data_b(1284) <= "0000000000";
data_b(1285) <= "0000000000";
data_b(1286) <= "0100000001";
data_b(1287) <= "0000000000";
data_b(1288) <= "0100000001";
data_b(1289) <= "0100000001";
data_b(1290) <= "0000000000";
data_b(1291) <= "0010000010";
data_b(1292) <= "0010000010";
data_b(1293) <= "0000000000";
data_b(1294) <= "0001000100";
data_b(1295) <= "0000000000";
--------------------------------81
data_b(1296) <= "0001000100";
data_b(1297) <= "0001000100";
data_b(1298) <= "0000000000";
data_b(1299) <= "0000000000";
data_b(1300) <= "0010000000";
data_b(1301) <= "0010000000";
data_b(1302) <= "0000000000";
data_b(1303) <= "0000000000";
data_b(1304) <= "1000000000";
data_b(1305) <= "1000000000";
data_b(1306) <= "0000000000";
data_b(1307) <= "0000000000";
data_b(1308) <= "0000000000";
data_b(1309) <= "0000000000";
data_b(1310) <= "0000000000";
data_b(1311) <= "0000000000";
-----------------------------------82
data_b(1312) <= "0001000010";
data_b(1313) <= "0001000010";
data_b(1314) <= "0000000000";
data_b(1315) <= "0000000000";
data_b(1316) <= "0000000000";
data_b(1317) <= "0000000000";
data_b(1318) <= "0010000100";
data_b(1319) <= "0010000100";
data_b(1320) <= "0000000000";
data_b(1321) <= "0000000000";
data_b(1322) <= "0000000000";
data_b(1323) <= "0000000000";
data_b(1324) <= "1000001000";
data_b(1325) <= "1000001000";
data_b(1326) <= "0000000000";
data_b(1327) <= "0000000000";
------------------------------83
data_b(1328) <= "0010001000";
data_b(1329) <= "0010001000";
data_b(1330) <= "0010000000";
data_b(1331) <= "0000000100";
data_b(1332) <= "0000000100";
data_b(1333) <= "0000000000";
data_b(1334) <= "0000001000";
data_b(1335) <= "0000000000";
data_b(1336) <= "0100001000";
data_b(1337) <= "0100001000";
data_b(1338) <= "0100000000";
data_b(1339) <= "0000000100";
data_b(1340) <= "0000000100";
data_b(1341) <= "0000000000";
data_b(1342) <= "0000001000";
data_b(1343) <= "0000000000";
------------------------------84
data_b(1344) <= "1000000100";
data_b(1345) <= "1000000100";
data_b(1346) <= "1000000100";
data_b(1347) <= "1000000100";
data_b(1348) <= "1000000100";
data_b(1349) <= "1000000100";
data_b(1350) <= "1000000100";
data_b(1351) <= "1000000100";
data_b(1352) <= "1000000100";
data_b(1353) <= "1000000100";
data_b(1354) <= "1000000100";
data_b(1355) <= "1000000100";
data_b(1356) <= "1000000100";
data_b(1357) <= "1000000100";
data_b(1358) <= "0000000000";
data_b(1359) <= "0000000000";
-----------------------------------85
----------------------------



		

process (n_clk,rss,rst)
begin
   if rss = '1' or rst = '1' then
      dot_data_00 <= zr;
		dot_data_01 <= zr;
		dot_data_02 <= zr;
		dot_data_03 <= zr;
		dot_data_04 <= zr;
		dot_data_05 <= zr;
		dot_data_06 <= zr;
		dot_data_07 <= zr;
		dot_data_08 <= zr;
		dot_data_09 <= zr;
		dot_data_10 <= zr;
		dot_data_11 <= zr;
		dot_data_12 <= zr;
		dot_data_13 <= zr;
		d_dp <= zr;
		d_d  <= zr;
		d_dm <= zr;
	elsif n_clk'event and n_clk = '1' then
		d_dp        <= dot_data_00;
		d_d         <= dot_data_01;
		d_dm        <= dot_data_02;
		dot_data_00 <= dot_data_01;
		dot_data_01 <= dot_data_02;
		dot_data_02 <= dot_data_03;
		dot_data_03 <= dot_data_04;
		dot_data_04 <= dot_data_05;
		dot_data_05 <= dot_data_06;
		dot_data_06 <= dot_data_07;
		dot_data_07 <= dot_data_08;
		dot_data_08 <= dot_data_09;
		dot_data_09 <= dot_data_10;
		dot_data_10 <= dot_data_11;
		dot_data_11 <= dot_data_12;
		dot_data_12 <= dot_data_13;
		dot_data_13 <= data_b(note);
	end if;
end process;




u0 : dot_dis
port map (
	clk => clk,
	dot_data_00 => dot_data_00,
	dot_data_01 => dot_data_01,
	dot_data_02 => dot_data_02,
	dot_data_03 => dot_data_03,
	dot_data_04 => dot_data_04,
	dot_data_05 => dot_data_05,
	dot_data_06 => dot_data_06,
	dot_data_07 => dot_data_07,
	dot_data_08 => dot_data_08,
	dot_data_09 => dot_data_09,
	dot_data_10 => dot_data_10,
	dot_data_11 => dot_data_11,
	dot_data_12 => dot_data_12,
	dot_data_13 => dot_data_13,
	dot_d => dot_d,
	dot_scan => dot_scan 
);

led <= st;



end a;