----------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

entity bubble_easy is
port (
	clk		: in std_logic;     -- 25MHz
	p1       : in std_logic;
	rss      : in std_logic;
	note_clk : out std_logic;
	d_d      : out std_logic_vector(9 downto 0);
	d_dp     : out std_logic_vector(9 downto 0);
	d_dm     : out std_logic_vector(9 downto 0);	
	reset    : out std_logic;	
	rr       : in std_logic;
   -------------------------------------------------------dot port
	dot_d : out std_logic_vector ( 9 downto 0);
	dot_scan : out std_logic_vector ( 13 downto 0);
	--------------------------------------------------------piezo port
	piezo	   : out std_logic;
	piezo2   : out std_logic;
	led : out std_logic
);
end bubble_easy;

----------------------------------------------------------------------------------
architecture a of bubble_easy is
-------------------------------------------------------------------------------component
component dot_dis
port (
	clk : in std_logic;
	dot_data_00 : in std_logic_vector (9 downto 0);
	dot_data_01 : in std_logic_vector (9 downto 0);
	dot_data_02 : in std_logic_vector (9 downto 0);
	dot_data_03 : in std_logic_vector (9 downto 0);
	dot_data_04 : in std_logic_vector (9 downto 0);
	dot_data_05 : in std_logic_vector (9 downto 0);
	dot_data_06 : in std_logic_vector (9 downto 0);
	dot_data_07 : in std_logic_vector (9 downto 0);
	dot_data_08 : in std_logic_vector (9 downto 0);
	dot_data_09 : in std_logic_vector (9 downto 0);
	dot_data_10 : in std_logic_vector (9 downto 0);
	dot_data_11 : in std_logic_vector (9 downto 0);
	dot_data_12 : in std_logic_vector (9 downto 0);
	dot_data_13 : in std_logic_vector (9 downto 0);

	dot_d : out std_logic_vector (9 downto 0);
	dot_scan : out std_logic_vector ( 13 downto 0)
);
end component;
------------------------------------------------------------------------com signal
signal ryt  : integer range 0 to 620312;
signal note : integer range 0 to 1700 := 1650;
signal n_clk   : std_logic := '0';
signal rst : std_logic := '0';

---------------------------------------------------------------------dot signal
signal dot_data_00 : std_logic_vector (9 downto 0);
signal dot_data_01 : std_logic_vector (9 downto 0);
signal dot_data_02 : std_logic_vector (9 downto 0);
signal dot_data_03 : std_logic_vector (9 downto 0);
signal dot_data_04 : std_logic_vector (9 downto 0);
signal dot_data_05 : std_logic_vector (9 downto 0);
signal dot_data_06 : std_logic_vector (9 downto 0);
signal dot_data_07 : std_logic_vector (9 downto 0);
signal dot_data_08 : std_logic_vector (9 downto 0);
signal dot_data_09 : std_logic_vector (9 downto 0);
signal dot_data_10 : std_logic_vector (9 downto 0);
signal dot_data_11 : std_logic_vector (9 downto 0);
signal dot_data_12 : std_logic_vector (9 downto 0);
signal dot_data_13 : std_logic_vector (9 downto 0);

constant zr : std_logic_vector(9 downto 0) := "0000000000";

type data_a is array(1700 downto 0) of std_logic_vector(9 downto 0);
signal data_b : data_a;

--------------------------------------------------------------------piezo signal
constant r  : integer range 0 to 1000000 := 0;

constant a_1 	: integer range 0 to 1000000 := 454544;
constant bm_1 	: integer range 0 to 1000000 := 429034;
constant b_1 	: integer range 0 to 1000000 := 404954;
constant c_1 	: integer range 0 to 1000000 := 382226;
constant dm_1 	: integer range 0 to 1000000 := 360773;
constant d_1 	: integer range 0 to 1000000 := 340524;
constant em_1 	: integer range 0 to 1000000 := 321414;
constant e_1 	: integer range 0 to 1000000 := 303373;
constant f_1 	: integer range 0 to 1000000 := 286346;
constant gm_1 	: integer range 0 to 1000000 := 270274;
constant g_1 	: integer range 0 to 1000000 := 255105;
constant am_1 	: integer range 0 to 1000000 := 240787;

constant a_2 	: integer range 0 to 1000000 := 227273;
constant bm_2 	: integer range 0 to 1000000 := 214517;
constant b_2 	: integer range 0 to 1000000 := 202477;
constant c_2 	: integer range 0 to 1000000 := 191113;
constant dm_2 	: integer range 0 to 1000000 := 180387;
constant d_2 	: integer range 0 to 1000000 := 170262;
constant em_2 	: integer range 0 to 1000000 := 160706;
constant e_2 	: integer range 0 to 1000000 := 151686;
constant f_2 	: integer range 0 to 1000000 := 143173;
constant gm_2 	: integer range 0 to 1000000 := 135137;
constant g_2 	: integer range 0 to 1000000 := 127553;
constant am_2 	: integer range 0 to 1000000 := 120394;

constant a_3 	: integer range 0 to 1000000 := 113635;
constant bm_3 	: integer range 0 to 1000000 := 107257;
constant b_3 	: integer range 0 to 1000000 := 101237;
constant c_3 	: integer range 0 to 1000000 := 95555;
constant dm_3 	: integer range 0 to 1000000 := 90192;
constant d_3 	: integer range 0 to 1000000 := 85130;
constant em_3 	: integer range 0 to 1000000 := 80352;
constant e_3 	: integer range 0 to 1000000 := 75842;
constant f_3 	: integer range 0 to 1000000 := 71585;
constant gm_3 	: integer range 0 to 1000000 := 67568;
constant g_3 	: integer range 0 to 1000000 := 63775;
constant am_3 	: integer range 0 to 1000000 := 60196;

constant a_4 	: integer range 0 to 1000000 := 56817;
constant bm_4 	: integer range 0 to 1000000 := 53628;
constant b_4 	: integer range 0 to 1000000 := 50618;
constant c_4 	: integer range 0 to 1000000 := 47777;
constant dm_4 	: integer range 0 to 1000000 := 45096;
constant d_4 	: integer range 0 to 1000000 := 42565;
constant em_4 	: integer range 0 to 1000000 := 40176;
constant e_4 	: integer range 0 to 1000000 := 37921;
constant f_4 	: integer range 0 to 1000000 := 35792;
constant gm_4 	: integer range 0 to 1000000 := 33783;
constant g_4 	: integer range 0 to 1000000 := 31887;
constant am_4 	: integer range 0 to 1000000 := 30097;

constant a_5 	: integer range 0 to 1000000 := 28408;
constant bm_5 	: integer range 0 to 1000000 := 26814;
constant b_5 	: integer range 0 to 1000000 := 25309;
constant c_5 	: integer range 0 to 1000000 := 23888;
constant dm_5 	: integer range 0 to 1000000 := 22547;
constant d_5 	: integer range 0 to 1000000 := 21282;
constant em_5 	: integer range 0 to 1000000 := 20087;
constant e_5 	: integer range 0 to 1000000 := 18960;
constant f_5 	: integer range 0 to 1000000 := 17896;
constant gm_5 	: integer range 0 to 1000000 := 16891;
constant g_5 	: integer range 0 to 1000000 := 15943;
constant am_5 	: integer range 0 to 1000000 := 15048;

constant a_6 	: integer range 0 to 1000000 := 14204;
constant bm_6 	: integer range 0 to 1000000 := 13406;
constant b_6 	: integer range 0 to 1000000 := 12654;
constant c_6 	: integer range 0 to 1000000 := 11945;
constant dm_6 	: integer range 0 to 1000000 := 11273;
constant d_6 	: integer range 0 to 1000000 := 10640;
constant em_6 	: integer range 0 to 1000000 := 10043;
constant e_6 	: integer range 0 to 1000000 := 9479;
constant f_6 	: integer range 0 to 1000000 := 8947;
constant gm_6 	: integer range 0 to 1000000 := 8445;
constant g_6 	: integer range 0 to 1000000 := 7971;
constant am_6 	: integer range 0 to 1000000 := 7524;


signal cnt 	: integer range 0 to 1000000;
signal cnt2 : integer range 0 to 1000000;
signal seq  : integer range 0 to 100000;


signal st   : std_logic := '0';

signal p_clk	: std_logic;
signal p_clk2  : std_logic;

type scale_a is array (1700 downto 0) of integer range 0 to 1000000;
signal scale : scale_a;
signal scale2: scale_a;
------------------------------------------------------------------------com

begin

process(p1,rss,rst)
begin
  if p1 = '1' then
     st <= '1';
  elsif rst = '1' or rss = '1' then
     st <= '0';
	  seq <= 0;
  end if;
end process;

process(clk,rst,rss)
begin
  if rst = '1' or rss = '1' then
     ryt <= 0;
	  n_clk <= '0';
  elsif clk'event and clk = '1' and st = '1' then
     if ryt = 620312 then
	     ryt <= 0;
        n_clk <= not n_clk;
     else
        ryt <= ryt + 1;
        n_clk <= n_clk;		  
     end if;
  end if;
end process;

note_clk <= n_clk;

process(n_clk,rss,rst,clk)
begin
  if rss = '1' or rst = '1' then
     note <= 1650;
  elsif n_clk'event and n_clk = '1' then
     if note = 1640 then
	     note <= 1650;
		  rst <= '1';
	  elsif note = 1700 then
	     note <= 0;
	  else
		  note <= note + 1;
     end if;
  end if;
  if rss = '1' or rr = '1' then
     rst <= '0';
  end if;  
end process;
reset <= rst;

---------------------------------------------------------------------dot
data_b(0) <= "0000000001";
data_b(1) <= "0000000000";
data_b(2) <= "0000000000";
data_b(3) <= "0000000000";
data_b(4) <= "0000000010";
data_b(5) <= "0000000000";
data_b(6) <= "0000000000";
data_b(7) <= "0000000000";
data_b(8) <= "0000000100";
data_b(9) <= "0000000100";
data_b(10) <= "0000000000";
data_b(11) <= "0000000000";
data_b(12) <= "0000000000";
data_b(13) <= "0000000000";
data_b(14) <= "0010000000";
data_b(15) <= "0000000000";
data_b(16) <= "0000000001";
data_b(17) <= "0000000000";
data_b(18) <= "0000000000";
data_b(19) <= "0000000000";
data_b(20) <= "0000000010";
data_b(21) <= "0000000000";
data_b(22) <= "0000000000";
data_b(23) <= "0000000000";
data_b(24) <= "0010000000";
data_b(25) <= "0000000000";
data_b(26) <= "0000000000";
data_b(27) <= "0000000000";
data_b(28) <= "0100000000";
data_b(29) <= "0000000000";
data_b(30) <= "0000000000";
data_b(31) <= "0000000000";
------------------------------------------------------------------------1����
data_b(32) <= "0000000001";
data_b(33) <= "0000000000";
data_b(34) <= "0000000000";
data_b(35) <= "0000000000";
data_b(36) <= "0000000010";
data_b(37) <= "0000000000";
data_b(38) <= "0000000000";
data_b(39) <= "0000000000";
data_b(40) <= "0000000100";
data_b(41) <= "0000000000";
data_b(42) <= "0010000000";
data_b(43) <= "0010000000";
data_b(44) <= "0000000000";
data_b(45) <= "0000000000";
data_b(46) <= "0000000000";
data_b(47) <= "0000000000";
data_b(48) <= "0000000010";
data_b(49) <= "0000000010";
data_b(50) <= "0000000010";
data_b(51) <= "0000000000";
data_b(52) <= "0000000000";
data_b(53) <= "0000000000";
data_b(54) <= "0000000000";
data_b(55) <= "0000000000";
data_b(56) <= "0000000000";
data_b(57) <= "0000000000";
data_b(58) <= "0000000000";
data_b(59) <= "0000000000";
data_b(60) <= "0000000100";
data_b(61) <= "0000000000";
data_b(62) <= "0010000000";
data_b(63) <= "0000000000";

------------------------------------------------------------------------2����
data_b(64) <= "1000000000";
data_b(65) <= "0000000000";
data_b(66) <= "0000000000";
data_b(67) <= "0000000000";
data_b(68) <= "0100000000";
data_b(69) <= "0000000000";
data_b(70) <= "0000000000";
data_b(71) <= "0000000000";
data_b(72) <= "0010000000";
data_b(73) <= "0000000000";
data_b(74) <= "0000000000";
data_b(75) <= "0000000000";
data_b(76) <= "0000000100";
data_b(77) <= "0000000000";
data_b(78) <= "0000000000";
data_b(79) <= "0000000000";
data_b(80) <= "0100000000";
data_b(81) <= "0000000000";
data_b(82) <= "0000000000";
data_b(83) <= "0000000000";
data_b(84) <= "0010000000";
data_b(85) <= "0000000000";
data_b(86) <= "0000000100";
data_b(87) <= "0000000100";
data_b(88) <= "0000000000";
data_b(89) <= "0000000000";
data_b(90) <= "0000000000";
data_b(91) <= "0000000000";
data_b(92) <= "0000000010";
data_b(93) <= "0000000000";
data_b(94) <= "0000000000";
data_b(95) <= "0000000000";
---------------------------------------------------------- 3����
data_b(96) <= "1000000000";
data_b(97) <= "0000000000";
data_b(98) <= "0000000000";
data_b(99) <= "0000000000";
data_b(100) <= "0100000000";
data_b(101) <= "0000000000";
data_b(102) <= "0000000000";
data_b(103) <= "0000000000";
data_b(104) <= "0010000000";
data_b(105) <= "0000000000";
data_b(106) <= "0100000000";
data_b(107) <= "0100000000";
data_b(108) <= "0000000000";
data_b(109) <= "0000000000";
data_b(110) <= "0000000000";
data_b(111) <= "0000000000";
data_b(112) <= "1000000000";
data_b(113) <= "0000000000";
data_b(114) <= "0000000000";
data_b(115) <= "0000000000";
data_b(116) <= "1000000000";
data_b(117) <= "0000000000";
data_b(118) <= "0000000000";
data_b(119) <= "0000000000";
data_b(120) <= "0100000000";
data_b(121) <= "0000000000";
data_b(122) <= "0000000000";
data_b(123) <= "0000000000";
data_b(124) <= "0010000000";
data_b(125) <= "0000000000";
data_b(126) <= "0000000000";
data_b(127) <= "0000000000";
-------------------------------------------------------------4����
data_b(128) <= "0000000100";
data_b(129) <= "0000000000";
data_b(130) <= "0000000000";
data_b(131) <= "0000000000";
data_b(132) <= "0010000000";
data_b(133) <= "0000000000";
data_b(134) <= "0000000000";
data_b(135) <= "0000000000";
data_b(136) <= "0100000000";
data_b(137) <= "0100000000";
data_b(138) <= "0000000000";
data_b(139) <= "0000000000";
data_b(140) <= "0000000000";
data_b(141) <= "0000000000";
data_b(142) <= "1000000000";
data_b(143) <= "0000000000";
data_b(144) <= "0000000001";
data_b(145) <= "0000000000";
data_b(146) <= "0000000000";
data_b(147) <= "0000000000";
data_b(148) <= "0000000010";
data_b(149) <= "0000000000";
data_b(150) <= "0000000000";
data_b(151) <= "0000000000";
data_b(152) <= "0000000100";
data_b(153) <= "0000000000";
data_b(154) <= "0010000000";
data_b(155) <= "0010000000";
data_b(156) <= "0000000000";
data_b(157) <= "0000000000";
data_b(158) <= "0000000000";
data_b(159) <= "0000000000";
------------------------------------------------------------------5����
data_b(160) <= "0000000001";
data_b(161) <= "0000000000";
data_b(162) <= "0000000000";
data_b(163) <= "0000000000";
data_b(164) <= "0000000010";
data_b(165) <= "0000000000";
data_b(166) <= "0000000000";
data_b(167) <= "0000000000";
data_b(168) <= "0000000100";
data_b(169) <= "0000000000";
data_b(170) <= "0010000000";
data_b(171) <= "0010000000";
data_b(172) <= "0000000000";
data_b(173) <= "0000000000";
data_b(174) <= "0000000000";
data_b(175) <= "0000000000";
data_b(176) <= "0000000010";
data_b(177) <= "0000000010";
data_b(178) <= "0000000010";
data_b(179) <= "0000000000";
data_b(180) <= "0000000000";
data_b(181) <= "0000000000";
data_b(182) <= "0000000000";
data_b(183) <= "0000000000";
data_b(184) <= "0000000000";
data_b(185) <= "0000000000";
data_b(186) <= "0000000000";
data_b(187) <= "0000000000";
data_b(188) <= "0000000100";
data_b(189) <= "0000000000";
data_b(190) <= "0010000000";
data_b(191) <= "0000000000";
----------------------------------------------------------------------6����
data_b(192) <= "1000000000";
data_b(193) <= "0000000000";
data_b(194) <= "0000000000";
data_b(195) <= "0000000000";
data_b(196) <= "0100000000";
data_b(197) <= "0000000000";
data_b(198) <= "0000000000";
data_b(199) <= "0000000000";
data_b(200) <= "0010000000";
data_b(201) <= "0000000000";
data_b(202) <= "0000000000";
data_b(203) <= "0000000000";
data_b(204) <= "0000000100";
data_b(205) <= "0000000000";
data_b(206) <= "0000000000";
data_b(207) <= "0000000000";
data_b(208) <= "0100000000";
data_b(209) <= "0000000000";
data_b(210) <= "0000000000";
data_b(211) <= "0000000000";
data_b(212) <= "0010000000";
data_b(213) <= "0000000000";
data_b(214) <= "0000000100";
data_b(215) <= "0000000100";
data_b(216) <= "0000000000";
data_b(217) <= "0000000000";
data_b(218) <= "0000000000";
data_b(219) <= "0000000000";
data_b(220) <= "0000000010";
data_b(221) <= "0000000000";
data_b(222) <= "0000000000";
data_b(223) <= "0000000000";
--------------------------------------------------7����
data_b(224) <= "1000000000";
data_b(225) <= "0000000000";
data_b(226) <= "0000000000";
data_b(227) <= "0000000000";
data_b(228) <= "0100000000";
data_b(229) <= "0000000000";
data_b(230) <= "0000000000";
data_b(231) <= "0000000000";
data_b(232) <= "0010000000";
data_b(233) <= "0000000000";
data_b(234) <= "1000000000";
data_b(235) <= "1000000000";
data_b(236) <= "0000000000";
data_b(237) <= "0000000000";
data_b(238) <= "0000000000";
data_b(239) <= "0000000000";
data_b(240) <= "0000000100";
data_b(241) <= "0000000000";
data_b(242) <= "0000000000";
data_b(243) <= "0000000000";
data_b(244) <= "1000000000";
data_b(245) <= "0000000000";
data_b(246) <= "0000000000";
data_b(247) <= "0000000000";
data_b(248) <= "0100000000";
data_b(249) <= "0000000000";
data_b(250) <= "0000000000";
data_b(251) <= "0000000000";
data_b(252) <= "0010000000";
data_b(253) <= "0000000000";
data_b(254) <= "0000000000";
data_b(255) <= "0000000000";
----------------------------------------------8����
data_b(256) <= "1000000000";          
data_b(257) <= "1000000000";
data_b(258) <= "1000000000";
data_b(259) <= "1000000000";
data_b(260) <= "1000000000";
data_b(261) <= "1000000000";
data_b(262) <= "1000000000";
data_b(263) <= "1000000000";
data_b(264) <= "1010000000";
data_b(265) <= "1000000000";
data_b(266) <= "1000000000";
data_b(267) <= "1000000000";
data_b(268) <= "1000000100";
data_b(269) <= "1000000000";
data_b(270) <= "1000000000";
data_b(271) <= "1000000000";
data_b(272) <= "0000000010";
data_b(273) <= "0000000000";
data_b(274) <= "0000000000";
data_b(275) <= "0000000000";
data_b(276) <= "0000000100";
data_b(277) <= "0000000000";
data_b(278) <= "0000000000";
data_b(279) <= "0000000000";
data_b(280) <= "0000000010";
data_b(281) <= "0000000000";
data_b(282) <= "0000000000";
data_b(283) <= "0000000000";
data_b(284) <= "0000000001";
data_b(285) <= "0000000000";
data_b(286) <= "0000000000";
data_b(287) <= "0000000000";
----------------------------------------------9����
data_b(288) <= "1000000000";          
data_b(289) <= "1000000000";
data_b(290) <= "1000000000";
data_b(291) <= "1000000000";
data_b(292) <= "1000000000";
data_b(293) <= "1000000000";
data_b(294) <= "1000000000";
data_b(295) <= "1000000000";
data_b(296) <= "1010000000";
data_b(297) <= "1000000000";
data_b(298) <= "1000000000";
data_b(299) <= "1000000000";
data_b(300) <= "1000000100";
data_b(301) <= "1000000000";
data_b(302) <= "1000000000";
data_b(303) <= "1000000000";
data_b(304) <= "0000000010";
data_b(305) <= "0000000000";
data_b(306) <= "0000000000";
data_b(307) <= "0000000000";
data_b(308) <= "0000000100";
data_b(309) <= "0000000000";
data_b(310) <= "0000000000";
data_b(311) <= "0000000000";
data_b(312) <= "0000000010";
data_b(313) <= "0000000000";
data_b(314) <= "0000000000";
data_b(315) <= "0000000000";
data_b(316) <= "0000000001";
data_b(317) <= "0000000000";
data_b(318) <= "0000000000";
data_b(319) <= "0000000000";
---------------------------------------------10����
data_b(320) <= "1000000000";          
data_b(321) <= "1000000000";
data_b(322) <= "1000000000";
data_b(323) <= "1000000000";
data_b(324) <= "1000000000";
data_b(325) <= "1000000000";
data_b(326) <= "1000000000";
data_b(327) <= "1000000000";
data_b(328) <= "1010000000";
data_b(329) <= "1000000000";
data_b(330) <= "1000000000";
data_b(331) <= "1000000000";
data_b(332) <= "1000000100";
data_b(333) <= "1000000000";
data_b(334) <= "1000000000";
data_b(335) <= "1000000000";
data_b(336) <= "0000000010";
data_b(337) <= "0000000000";
data_b(338) <= "0000000000";
data_b(339) <= "0000000000";
data_b(340) <= "0000000100";
data_b(341) <= "0000000000";
data_b(342) <= "0000000000";
data_b(343) <= "0000000000";
data_b(344) <= "0000000010";
data_b(345) <= "0000000000";
data_b(346) <= "0000000000";
data_b(347) <= "0000000000";
data_b(348) <= "0000000001";
data_b(349) <= "0000000000";
data_b(350) <= "0000000000";
data_b(351) <= "0000000000";
-----------------------------------------------11����
data_b(352) <= "1000000000";          
data_b(353) <= "1000000000";
data_b(354) <= "1000000000";
data_b(355) <= "1000000000";
data_b(356) <= "1000000000";
data_b(357) <= "1000000000";
data_b(358) <= "1000000000";
data_b(359) <= "1000000000";
data_b(360) <= "1010000000";
data_b(361) <= "1000000000";
data_b(362) <= "1000000000";
data_b(363) <= "1000000000";
data_b(364) <= "1000000100";
data_b(365) <= "1000000000";
data_b(366) <= "1000000000";
data_b(367) <= "1000000000";
data_b(368) <= "0000000010";
data_b(369) <= "0000000000";
data_b(370) <= "0000000000";
data_b(371) <= "0000000000";
data_b(372) <= "0000000100";
data_b(373) <= "0000000000";
data_b(374) <= "0000000000";
data_b(375) <= "0000000000";
data_b(376) <= "0000000010";
data_b(377) <= "0000000000";
data_b(378) <= "0000000000";
data_b(379) <= "0000000000";
data_b(380) <= "0000000001";
data_b(381) <= "0000000000";
data_b(382) <= "0000000000";
data_b(383) <= "0000000000";
-----------------------------------------------12����
data_b(384) <= "0000000001";
data_b(385) <= "0000000000";
data_b(386) <= "0000000000";
data_b(387) <= "0000000000";
data_b(388) <= "0000000001";
data_b(389) <= "0000000001";
data_b(390) <= "0000000000";
data_b(391) <= "0000000000";
data_b(392) <= "0000000000";
data_b(393) <= "0000000000";
data_b(394) <= "0000000000";
data_b(395) <= "0000000000";
data_b(396) <= "0000000001";
data_b(397) <= "0000000001";
data_b(398) <= "0000000000";
data_b(399) <= "0000000000";
data_b(400) <= "0000000000";
data_b(401) <= "0000000000";
data_b(402) <= "0000000000";
data_b(403) <= "0000000000";
data_b(404) <= "0000000010";
data_b(405) <= "0000000000";
data_b(406) <= "0000000000";
data_b(407) <= "0000000000";
data_b(408) <= "0000000100";
data_b(409) <= "0000000100";
data_b(410) <= "0000000000";
data_b(411) <= "0000000000";
data_b(412) <= "0000000000";
data_b(413) <= "0000000000";
data_b(414) <= "0000000000";
data_b(415) <= "0000000000";
------------------------------------------------------13����
data_b(416) <= "0000000010";
data_b(417) <= "0000000010";
data_b(418) <= "0000000010";
data_b(419) <= "0000000010";
data_b(420) <= "0000000010";
data_b(421) <= "0000000010";
data_b(422) <= "0000000010";
data_b(423) <= "0000000010";
data_b(424) <= "0000000010";
data_b(425) <= "0000000010";
data_b(426) <= "0000000010";
data_b(427) <= "0000000010";
data_b(428) <= "0000000000";
data_b(429) <= "0000000000";
data_b(430) <= "0000000000";
data_b(431) <= "0000000000";
data_b(432) <= "0000000000";
data_b(433) <= "0000000000";
data_b(434) <= "0000000000";
data_b(435) <= "0000000000";
data_b(436) <= "0000000000";
data_b(437) <= "0000000000";
data_b(438) <= "0000000000";
data_b(439) <= "0000000000";
data_b(440) <= "0000000010";
data_b(441) <= "0000000010";
data_b(442) <= "0000000010";
data_b(443) <= "0000000010";
data_b(444) <= "0000000000";
data_b(445) <= "0000000000";
data_b(446) <= "0000000000";
data_b(447) <= "0000000000";
-------------------------------------------------------14����
data_b(448) <= "0000000100";
data_b(449) <= "0000000100";
data_b(450) <= "0000000100";
data_b(451) <= "0000000000";
data_b(452) <= "0000000000";
data_b(453) <= "0000000000";
data_b(454) <= "0000000000";
data_b(455) <= "0000000000";
data_b(456) <= "0000000000";
data_b(457) <= "0000000000";
data_b(458) <= "0000000000";
data_b(459) <= "0000000000";
data_b(460) <= "1000000000";
data_b(461) <= "1000000000";
data_b(462) <= "0000000000";
data_b(463) <= "0000000000";
data_b(464) <= "0000000000";
data_b(465) <= "0000000000";
data_b(466) <= "0000000000";
data_b(467) <= "0000000000";
data_b(468) <= "1000000000";
data_b(469) <= "0000000000";
data_b(470) <= "0000000000";
data_b(471) <= "0000000000";
data_b(472) <= "0000000010";
data_b(473) <= "0000000010";
data_b(474) <= "0000000000";
data_b(475) <= "0000000000";
data_b(476) <= "0000000000";
data_b(477) <= "0000000000";
data_b(478) <= "0000000000";
data_b(479) <= "0000000000";
------------------------------------------------------15����
data_b(480) <= "0000000010";                                   
data_b(481) <= "0000000010";
data_b(482) <= "0000000010";
data_b(483) <= "0000000010";
data_b(484) <= "0000000010";
data_b(485) <= "0000000010";
data_b(486) <= "0000000010";
data_b(487) <= "0000000010";
data_b(488) <= "0000000010";
data_b(489) <= "0000000010";
data_b(490) <= "0000000000";
data_b(491) <= "0000000000";
data_b(492) <= "0000000000";
data_b(493) <= "0000000000";
data_b(494) <= "0000000000";
data_b(495) <= "0000000000";
data_b(496) <= "0000000000";
data_b(497) <= "0000000000";
data_b(498) <= "0000000000";
data_b(499) <= "0000000000";
data_b(500) <= "1000000000";
data_b(501) <= "0000000000";
data_b(502) <= "0000000000";
data_b(503) <= "0000000000";
data_b(504) <= "0100000000";
data_b(505) <= "0000000000";
data_b(506) <= "0000000000";
data_b(507) <= "0000000000";
data_b(508) <= "0010000000";
data_b(509) <= "0000000000";
data_b(510) <= "0000000000";
data_b(511) <= "0000000000";
-------------------------------------------------------16����
data_b(512) <= "1000000000";          
data_b(513) <= "1000000000";
data_b(514) <= "1000000000";
data_b(515) <= "1000000000";
data_b(516) <= "1000000000";
data_b(517) <= "1000000000";
data_b(518) <= "1000000000";
data_b(519) <= "1000000000";
data_b(520) <= "1010000000";
data_b(521) <= "1000000000";
data_b(522) <= "1000000000";
data_b(523) <= "1000000000";
data_b(524) <= "1000000100";
data_b(525) <= "1000000000";
data_b(526) <= "1000000000";
data_b(527) <= "1000000000";
data_b(528) <= "0000000010";
data_b(529) <= "0000000000";
data_b(530) <= "0000000000";
data_b(531) <= "0000000000";
data_b(532) <= "0000000100";
data_b(533) <= "0000000000";
data_b(534) <= "0000000000";
data_b(535) <= "0000000000";
data_b(536) <= "0000000010";
data_b(537) <= "0000000000";
data_b(538) <= "0000000000";
data_b(539) <= "0000000000";
data_b(540) <= "0000000001";
data_b(541) <= "0000000000";
data_b(542) <= "0000000000";
data_b(543) <= "0000000000";
---------------------------------------------------------17����
data_b(544) <= "1000000000";          
data_b(545) <= "1000000000";
data_b(546) <= "1000000000";
data_b(547) <= "1000000000";
data_b(548) <= "1000000000";
data_b(549) <= "1000000000";
data_b(550) <= "1000000000";
data_b(551) <= "1000000000";
data_b(552) <= "1010000000";
data_b(553) <= "1000000000";
data_b(554) <= "1000000000";
data_b(555) <= "1000000000";
data_b(556) <= "1000000100";
data_b(557) <= "1000000000";
data_b(558) <= "1000000000";
data_b(559) <= "1000000000";
data_b(560) <= "0000000010";
data_b(561) <= "0000000000";
data_b(562) <= "0000000000";
data_b(563) <= "0000000000";
data_b(564) <= "0000000100";
data_b(565) <= "0000000000";
data_b(566) <= "0000000000";
data_b(567) <= "0000000000";
data_b(568) <= "0000000010";
data_b(569) <= "0000000000";
data_b(570) <= "0000000000";
data_b(571) <= "0000000000";
data_b(572) <= "0000000001";
data_b(573) <= "0000000000";
data_b(574) <= "0000000000";
data_b(575) <= "0000000000";
------------------------------------18����
data_b(576) <= "1000000000";          
data_b(577) <= "1000000000";
data_b(578) <= "1000000000";
data_b(579) <= "1000000000";
data_b(580) <= "1000000000";
data_b(581) <= "1000000000";
data_b(582) <= "1000000000";
data_b(583) <= "1000000000";
data_b(584) <= "1010000000";
data_b(585) <= "1000000000";
data_b(586) <= "1000000000";
data_b(587) <= "1000000000";
data_b(588) <= "1000000100";
data_b(589) <= "1000000000";
data_b(590) <= "1000000000";
data_b(591) <= "1000000000";
data_b(592) <= "0000000010";
data_b(593) <= "0000000000";
data_b(594) <= "0000000000";
data_b(595) <= "0000000000";
data_b(596) <= "0000000100";
data_b(597) <= "0000000000";
data_b(598) <= "0000000000";
data_b(599) <= "0000000000";
data_b(600) <= "0000000010";
data_b(601) <= "0000000000";
data_b(602) <= "0000000000";
data_b(603) <= "0000000000";
data_b(604) <= "0000000001";
data_b(605) <= "0000000000";
data_b(606) <= "0000000000";
data_b(607) <= "0000000000";
------------------------------------------------------------19����
data_b(608) <= "1000000000";          
data_b(609) <= "1000000000";
data_b(610) <= "1000000000";
data_b(611) <= "1000000000";
data_b(612) <= "1000000000";
data_b(613) <= "1000000000";
data_b(614) <= "1000000000";
data_b(615) <= "1000000000";
data_b(616) <= "1010000000";
data_b(617) <= "1000000000";
data_b(618) <= "1000000000";
data_b(619) <= "1000000000";
data_b(620) <= "1000000100";
data_b(621) <= "1000000000";
data_b(622) <= "1000000000";
data_b(623) <= "1000000000";
data_b(624) <= "0000000010";
data_b(625) <= "0000000000";
data_b(626) <= "0000000000";
data_b(627) <= "0000000000";
data_b(628) <= "0000000100";
data_b(629) <= "0000000000";
data_b(630) <= "0000000000";
data_b(631) <= "0000000000";
data_b(632) <= "0000000010";
data_b(633) <= "0000000000";
data_b(634) <= "0000000000";
data_b(635) <= "0000000000";
data_b(636) <= "0000000001";
data_b(637) <= "0000000000";
data_b(638) <= "0000000000";
data_b(639) <= "0000000000";
------------------------------------------------------------------20����
data_b(640) <= "0000000001";
data_b(641) <= "0000000000";
data_b(642) <= "0000000000";
data_b(643) <= "0000000000";
data_b(644) <= "0000000001";
data_b(645) <= "0000000001";
data_b(646) <= "0000000000";
data_b(647) <= "0000000000";
data_b(648) <= "0000000000";
data_b(649) <= "0000000000";
data_b(650) <= "0000000000";
data_b(651) <= "0000000000";
data_b(652) <= "0000000001";
data_b(653) <= "0000000001";
data_b(654) <= "0000000000";
data_b(655) <= "0000000000";
data_b(656) <= "0000000000";
data_b(657) <= "0000000000";
data_b(658) <= "0000000000";
data_b(659) <= "0000000000";
data_b(660) <= "0000000010";
data_b(661) <= "0000000000";
data_b(662) <= "0000000000";
data_b(663) <= "0000000000";
data_b(664) <= "0000000100";
data_b(665) <= "0000000100";
data_b(666) <= "0000000000";
data_b(667) <= "0000000000";
data_b(668) <= "0000000000";
data_b(669) <= "0000000000";
data_b(670) <= "0000000000";
data_b(671) <= "0000000000";
------------------------------------21����

data_b(672) <= "0000000001";
data_b(673) <= "0000000001";
data_b(674) <= "0000000001";
data_b(675) <= "0000000001";
data_b(676) <= "0000000001";
data_b(677) <= "0000000001";
data_b(678) <= "0000000001";
data_b(679) <= "0000000001";
data_b(680) <= "0000000001";
data_b(681) <= "0000000001";
data_b(682) <= "0000000001";
data_b(683) <= "0000000001";
data_b(684) <= "0000000000";
data_b(685) <= "0000000000";
data_b(686) <= "0000000000";
data_b(687) <= "0000000000";
data_b(688) <= "0000000000";
data_b(689) <= "0000000000";
data_b(690) <= "0000000000";
data_b(691) <= "0000000000";
data_b(692) <= "0000000000";
data_b(693) <= "0000000000";
data_b(694) <= "0000000000";
data_b(695) <= "0000000000";
data_b(696) <= "0000000001";
data_b(697) <= "0000000001";
data_b(698) <= "0000000000";
data_b(699) <= "0000000000";
data_b(700) <= "0000000000";
data_b(701) <= "0000000000";
data_b(702) <= "0000000000";
data_b(703) <= "0000000000";
-----------------------------------------------------------22����
data_b(704) <= "0000000010";
data_b(705) <= "0000000010";
data_b(706) <= "0000000010";
data_b(707) <= "0000000000";
data_b(708) <= "0000000000";
data_b(709) <= "0000000000";
data_b(710) <= "0000000000";
data_b(711) <= "0000000000";
data_b(712) <= "0000000000";
data_b(713) <= "0000000000";
data_b(714) <= "0000000000";
data_b(715) <= "0000000000";
data_b(716) <= "1000000000";
data_b(717) <= "1000000000";
data_b(718) <= "0000000000";
data_b(719) <= "0000000000";
data_b(720) <= "0000000000";
data_b(721) <= "0000000000";
data_b(722) <= "0000000000";
data_b(723) <= "0000000000";
data_b(724) <= "0000000001";
data_b(725) <= "0000000000";
data_b(726) <= "0000000000";
data_b(727) <= "0000000000";
data_b(728) <= "1000000000";
data_b(729) <= "0000000000";
data_b(730) <= "0000000000";
data_b(731) <= "0000000000";
data_b(732) <= "0000000001";
data_b(733) <= "0000000000";
data_b(734) <= "0000000000";
data_b(735) <= "0000000000";
-----------------------------------------------------------------23����
data_b(736) <= "0000000100";
data_b(737) <= "0000000100";
data_b(738) <= "0000000100";
data_b(739) <= "0000000100";
data_b(740) <= "0000000100";
data_b(741) <= "0000000100";
data_b(742) <= "0000000100";
data_b(743) <= "0000000100";
data_b(744) <= "0000000100";
data_b(745) <= "0000000100";
data_b(746) <= "0000000000";
data_b(747) <= "0000000000";
data_b(748) <= "0000000000";
data_b(749) <= "0000000000";
data_b(750) <= "0000000000";
data_b(751) <= "0000000000";
data_b(752) <= "0000000000";
data_b(753) <= "0000000000";
data_b(754) <= "0000000000";
data_b(755) <= "0000000000";
data_b(756) <= "1000000000";
data_b(757) <= "0000000000";
data_b(758) <= "0000000000";
data_b(759) <= "0000000000";
data_b(760) <= "0100000000";
data_b(761) <= "0000000000";
data_b(762) <= "0000000000";
data_b(763) <= "0000000000";
data_b(764) <= "0010000000";
data_b(765) <= "0000000000";
data_b(766) <= "0000000000";
data_b(767) <= "0000000000";
---------------------------------------24����

---------------------------------------------------------------------dot
data_b(768) <= "0000000001";
data_b(769) <= "0000000000";
data_b(770) <= "0000000000";
data_b(771) <= "0000000000";
data_b(772) <= "0000000010";
data_b(773) <= "0000000000";
data_b(774) <= "0000000000";
data_b(775) <= "0000000000";
data_b(776) <= "0000000100";
data_b(777) <= "0000000100";
data_b(778) <= "0000000000";
data_b(779) <= "0000000000";
data_b(780) <= "0000000000";
data_b(781) <= "0000000000";
data_b(782) <= "0010000000";
data_b(783) <= "0000000000";
data_b(784) <= "0000000001";
data_b(785) <= "0000000000";
data_b(786) <= "0000000000";
data_b(787) <= "0000000000";
data_b(788) <= "0000000010";
data_b(789) <= "0000000000";
data_b(790) <= "0000000000";
data_b(791) <= "0000000000";
data_b(792) <= "0010000000";
data_b(793) <= "0000000000";
data_b(794) <= "0000000000";
data_b(795) <= "0000000000";
data_b(796) <= "0100000000";
data_b(797) <= "0000000000";
data_b(798) <= "0000000000";
data_b(799) <= "0000000000";
------------------------------------------------------------------------1����
data_b(800) <= "0000000001";
data_b(801) <= "0000000000";
data_b(802) <= "0000000000";
data_b(803) <= "0000000000";
data_b(804) <= "0000000010";
data_b(805) <= "0000000000";
data_b(806) <= "0000000000";
data_b(807) <= "0000000000";
data_b(808) <= "0000000100";
data_b(809) <= "0000000000";
data_b(810) <= "0010000000";
data_b(811) <= "0010000000";
data_b(812) <= "0000000000";
data_b(813) <= "0000000000";
data_b(814) <= "0000000000";
data_b(815) <= "0000000000";
data_b(816) <= "0000000010";
data_b(817) <= "0000000010";
data_b(818) <= "0000000010";
data_b(819) <= "0000000000";
data_b(820) <= "0000000000";
data_b(821) <= "0000000000";
data_b(822) <= "0000000000";
data_b(823) <= "0000000000";
data_b(824) <= "0000000000";
data_b(825) <= "0000000000";
data_b(826) <= "0000000000";
data_b(827) <= "0000000000";
data_b(828) <= "0000000100";
data_b(829) <= "0000000000";
data_b(830) <= "0010000000";
data_b(831) <= "0000000000";

------------------------------------------------------------------------2����
data_b(832) <= "1000000000";
data_b(833) <= "0000000000";
data_b(834) <= "0000000000";
data_b(835) <= "0000000000";
data_b(836) <= "0100000000";
data_b(837) <= "0000000000";
data_b(838) <= "0000000000";
data_b(839) <= "0000000000";
data_b(840) <= "0010000000";
data_b(841) <= "0000000000";
data_b(842) <= "0000000000";
data_b(843) <= "0000000000";
data_b(844) <= "0000000100";
data_b(845) <= "0000000000";
data_b(846) <= "0000000000";
data_b(847) <= "0000000000";
data_b(848) <= "0100000000";
data_b(849) <= "0000000000";
data_b(850) <= "0000000000";
data_b(851) <= "0000000000";
data_b(852) <= "0010000000";
data_b(853) <= "0000000000";
data_b(854) <= "0000000100";
data_b(855) <= "0000000100";
data_b(856) <= "0000000000";
data_b(857) <= "0000000000";
data_b(858) <= "0000000000";
data_b(859) <= "0000000000";
data_b(860) <= "0000000010";
data_b(861) <= "0000000000";
data_b(862) <= "0000000000";
data_b(863) <= "0000000000";
---------------------------------------------------------- 3����
data_b(864) <= "1000000000";
data_b(865) <= "0000000000";
data_b(866) <= "0000000000";
data_b(867) <= "0000000000";
data_b(868) <= "0100000000";
data_b(869) <= "0000000000";
data_b(870) <= "0000000000";
data_b(871) <= "0000000000";
data_b(872) <= "0010000000";
data_b(873) <= "0000000000";
data_b(874) <= "0100000000";
data_b(875) <= "0100000000";
data_b(876) <= "0000000000";
data_b(877) <= "0000000000";
data_b(878) <= "0000000000";
data_b(879) <= "0000000000";
data_b(880) <= "1000000000";
data_b(881) <= "0000000000";
data_b(882) <= "0000000000";
data_b(883) <= "0000000000";
data_b(884) <= "1000000000";
data_b(885) <= "0000000000";
data_b(886) <= "0000000000";
data_b(887) <= "0000000000";
data_b(888) <= "0100000000";
data_b(889) <= "0000000000";
data_b(890) <= "0000000000";
data_b(891) <= "0000000000";
data_b(892) <= "0010000000";
data_b(893) <= "0000000000";
data_b(894) <= "0000000000";
data_b(895) <= "0000000000";
-------------------------------------------------------------4����
data_b(896) <= "0000000100";
data_b(897) <= "0000000000";
data_b(898) <= "0000000000";
data_b(899) <= "0000000000";
data_b(900) <= "0010000000";
data_b(901) <= "0000000000";
data_b(902) <= "0000000000";
data_b(903) <= "0000000000";
data_b(904) <= "0100000000";
data_b(905) <= "0100000000";
data_b(906) <= "0000000000";
data_b(907) <= "0000000000";
data_b(908) <= "0000000000";
data_b(909) <= "0000000000";
data_b(910) <= "1000000000";
data_b(911) <= "0000000000";
data_b(912) <= "0000000001";
data_b(913) <= "0000000000";
data_b(914) <= "0000000000";
data_b(915) <= "0000000000";
data_b(916) <= "0000000010";
data_b(917) <= "0000000000";
data_b(918) <= "0000000000";
data_b(919) <= "0000000000";
data_b(920) <= "0000000100";
data_b(921) <= "0000000000";
data_b(922) <= "0010000000";
data_b(923) <= "0010000000";
data_b(924) <= "0000000000";
data_b(925) <= "0000000000";
data_b(926) <= "0000000000";
data_b(927) <= "0000000000";
------------------------------------------------------------------5����
data_b(928) <= "0000000001";
data_b(929) <= "0000000000";
data_b(930) <= "0000000000";
data_b(931) <= "0000000000";
data_b(932) <= "0000000010";
data_b(933) <= "0000000000";
data_b(934) <= "0000000000";
data_b(935) <= "0000000000";
data_b(936) <= "0000000100";
data_b(937) <= "0000000000";
data_b(938) <= "0010000000";
data_b(939) <= "0010000000";
data_b(940) <= "0000000000";
data_b(941) <= "0000000000";
data_b(942) <= "0000000000";
data_b(943) <= "0000000000";
data_b(944) <= "0000000010";
data_b(945) <= "0000000010";
data_b(946) <= "0000000010";
data_b(947) <= "0000000000";
data_b(948) <= "0000000000";
data_b(949) <= "0000000000";
data_b(950) <= "0000000000";
data_b(951) <= "0000000000";
data_b(952) <= "0000000000";
data_b(953) <= "0000000000";
data_b(954) <= "0000000000";
data_b(955) <= "0000000000";
data_b(956) <= "0000000100";
data_b(957) <= "0000000000";
data_b(958) <= "0010000000";
data_b(959) <= "0000000000";
----------------------------------------------------------------------6����
data_b(960) <= "1000000000";
data_b(961) <= "0000000000";
data_b(962) <= "0000000000";
data_b(963) <= "0000000000";
data_b(964) <= "0100000000";
data_b(965) <= "0000000000";
data_b(966) <= "0000000000";
data_b(967) <= "0000000000";
data_b(968) <= "0010000000";
data_b(969) <= "0000000000";
data_b(970) <= "0000000000";
data_b(971) <= "0000000000";
data_b(972) <= "0000000100";
data_b(973) <= "0000000000";
data_b(974) <= "0000000000";
data_b(975) <= "0000000000";
data_b(976) <= "0100000000";
data_b(977) <= "0000000000";
data_b(978) <= "0000000000";
data_b(979) <= "0000000000";
data_b(980) <= "0010000000";
data_b(981) <= "0000000000";
data_b(982) <= "0000000100";
data_b(983) <= "0000000100";
data_b(984) <= "0000000000";
data_b(985) <= "0000000000";
data_b(986) <= "0000000000";
data_b(987) <= "0000000000";
data_b(988) <= "0000000010";
data_b(989) <= "0000000000";
data_b(990) <= "0000000000";
data_b(991) <= "0000000000";
--------------------------------------------------7����
data_b(992) <= "1000000000";
data_b(993) <= "0000000000";
data_b(994) <= "0000000000";
data_b(995) <= "0000000000";
data_b(996) <= "0100000000";
data_b(997) <= "0000000000";
data_b(998) <= "0000000000";
data_b(999) <= "0000000000";
data_b(1000) <= "0010000000";
data_b(1001) <= "0000000000";
data_b(1002) <= "1000000000";
data_b(1003) <= "1000000000";
data_b(1004) <= "0000000000";
data_b(1005) <= "0000000000";
data_b(1006) <= "0000000000";
data_b(1007) <= "0000000000";
data_b(1008) <= "0000000100";
data_b(1009) <= "0000000000";
data_b(1010) <= "0000000000";
data_b(1011) <= "0000000000";
data_b(1012) <= "1000000000";
data_b(1013) <= "0000000000";
data_b(1014) <= "0000000000";
data_b(1015) <= "0000000000";
data_b(1016) <= "0100000000";
data_b(1017) <= "0000000000";
data_b(1018) <= "0000000000";
data_b(1019) <= "0000000000";
data_b(1020) <= "0010000000";
data_b(1021) <= "0000000000";
data_b(1022) <= "0000000000";
data_b(1023) <= "0000000000";
----------------------------------------------8����
data_b(1024) <= "1000000000";          
data_b(1025) <= "1000000000";
data_b(1026) <= "1000000000";
data_b(1027) <= "1000000000";
data_b(1028) <= "1000000000";
data_b(1029) <= "1000000000";
data_b(1030) <= "1000000000";
data_b(1031) <= "1000000000";
data_b(1032) <= "1010000000";
data_b(1033) <= "1000000000";
data_b(1034) <= "1000000000";
data_b(1035) <= "1000000000";
data_b(1036) <= "1000000100";
data_b(1037) <= "1000000000";
data_b(1038) <= "1000000000";
data_b(1039) <= "1000000000";
data_b(1040) <= "0000000010";
data_b(1041) <= "0000000000";
data_b(1042) <= "0000000000";
data_b(1043) <= "0000000000";
data_b(1044) <= "0000000100";
data_b(1045) <= "0000000000";
data_b(1046) <= "0000000000";
data_b(1047) <= "0000000000";
data_b(1048) <= "0000000010";
data_b(1049) <= "0000000000";
data_b(1050) <= "0000000000";
data_b(1051) <= "0000000000";
data_b(1052) <= "0000000001";
data_b(1053) <= "0000000000";
data_b(1054) <= "0000000000";
data_b(1055) <= "0000000000";
----------------------------------------------9����
data_b(1056) <= "1000000000";          
data_b(1057) <= "1000000000";
data_b(1058) <= "1000000000";
data_b(1059) <= "1000000000";
data_b(1060) <= "1000000000";
data_b(1061) <= "1000000000";
data_b(1062) <= "1000000000";
data_b(1063) <= "1000000000";
data_b(1064) <= "1010000000";
data_b(1065) <= "1000000000";
data_b(1066) <= "1000000000";
data_b(1067) <= "1000000000";
data_b(1068) <= "1000000100";
data_b(1069) <= "1000000000";
data_b(1070) <= "1000000000";
data_b(1071) <= "1000000000";
data_b(1072) <= "0000000010";
data_b(1073) <= "0000000000";
data_b(1074) <= "0000000000";
data_b(1075) <= "0000000000";
data_b(1076) <= "0000000100";
data_b(1077) <= "0000000000";
data_b(1078) <= "0000000000";
data_b(1079) <= "0000000000";
data_b(1080) <= "0000000010";
data_b(1081) <= "0000000000";
data_b(1082) <= "0000000000";
data_b(1083) <= "0000000000";
data_b(1084) <= "0000000001";
data_b(1085) <= "0000000000";
data_b(1086) <= "0000000000";
data_b(1087) <= "0000000000";
---------------------------------------------10����
data_b(1088) <= "1000000000";          
data_b(1089) <= "1000000000";
data_b(1090) <= "1000000000";
data_b(1091) <= "1000000000";
data_b(1092) <= "1000000000";
data_b(1093) <= "1000000000";
data_b(1094) <= "1000000000";
data_b(1095) <= "1000000000";
data_b(1096) <= "1010000000";
data_b(1097) <= "1000000000";
data_b(1098) <= "1000000000";
data_b(1099) <= "1000000000";
data_b(1100) <= "1000000100";
data_b(1101) <= "1000000000";
data_b(1102) <= "1000000000";
data_b(1103) <= "1000000000";
data_b(1104) <= "0000000010";
data_b(1105) <= "0000000000";
data_b(1106) <= "0000000000";
data_b(1107) <= "0000000000";
data_b(1108) <= "0000000100";
data_b(1109) <= "0000000000";
data_b(1110) <= "0000000000";
data_b(1111) <= "0000000000";
data_b(1112) <= "0000000010";
data_b(1113) <= "0000000000";
data_b(1114) <= "0000000000";
data_b(1115) <= "0000000000";
data_b(1116) <= "0000000001";
data_b(1117) <= "0000000000";
data_b(1118) <= "0000000000";
data_b(1119) <= "0000000000";
-----------------------------------------------11����
data_b(1120) <= "1000000000";          
data_b(1121) <= "1000000000";
data_b(1122) <= "1000000000";
data_b(1123) <= "1000000000";
data_b(1124) <= "1000000000";
data_b(1125) <= "1000000000";
data_b(1126) <= "1000000000";
data_b(1127) <= "1000000000";
data_b(1128) <= "1010000000";
data_b(1129) <= "1000000000";
data_b(1130) <= "1000000000";
data_b(1131) <= "1000000000";
data_b(1132) <= "1000000100";
data_b(1133) <= "1000000000";
data_b(1134) <= "1000000000";
data_b(1135) <= "1000000000";
data_b(1136) <= "0000000010";
data_b(1137) <= "0000000000";
data_b(1138) <= "0000000000";
data_b(1139) <= "0000000000";
data_b(1140) <= "0000000100";
data_b(1141) <= "0000000000";
data_b(1142) <= "0000000000";
data_b(1143) <= "0000000000";
data_b(1144) <= "0000000010";
data_b(1145) <= "0000000000";
data_b(1146) <= "0000000000";
data_b(1147) <= "0000000000";
data_b(1148) <= "0000000001";
data_b(1149) <= "0000000000";
data_b(1150) <= "0000000000";
data_b(1151) <= "0000000000";
-----------------------------------------------12����
data_b(1152) <= "0000000001";
data_b(1153) <= "0000000000";
data_b(1154) <= "0000000000";
data_b(1155) <= "0000000000";
data_b(1156) <= "0000000001";
data_b(1157) <= "0000000001";
data_b(1158) <= "0000000000";
data_b(1159) <= "0000000000";
data_b(1160) <= "0000000000";
data_b(1161) <= "0000000000";
data_b(1162) <= "0000000000";
data_b(1163) <= "0000000000";
data_b(1164) <= "0000000001";
data_b(1165) <= "0000000001";
data_b(1166) <= "0000000000";
data_b(1167) <= "0000000000";
data_b(1168) <= "0000000000";
data_b(1169) <= "0000000000";
data_b(1170) <= "0000000000";
data_b(1171) <= "0000000000";
data_b(1172) <= "0000000010";
data_b(1173) <= "0000000000";
data_b(1174) <= "0000000000";
data_b(1175) <= "0000000000";
data_b(1176) <= "0000000100";
data_b(1177) <= "0000000100";
data_b(1178) <= "0000000000";
data_b(1179) <= "0000000000";
data_b(1180) <= "0000000000";
data_b(1181) <= "0000000000";
data_b(1182) <= "0000000000";
data_b(1183) <= "0000000000";
------------------------------------------------------13����
data_b(1184) <= "0000000010";
data_b(1185) <= "0000000010";
data_b(1186) <= "0000000010";
data_b(1187) <= "0000000010";
data_b(1188) <= "0000000010";
data_b(1189) <= "0000000010";
data_b(1190) <= "0000000010";
data_b(1191) <= "0000000010";
data_b(1192) <= "0000000010";
data_b(1193) <= "0000000010";
data_b(1194) <= "0000000010";
data_b(1195) <= "0000000010";
data_b(1196) <= "0000000000";
data_b(1197) <= "0000000000";
data_b(1198) <= "0000000000";
data_b(1199) <= "0000000000";
data_b(1200) <= "0000000000";
data_b(1201) <= "0000000000";
data_b(1202) <= "0000000000";
data_b(1203) <= "0000000000";
data_b(1204) <= "0000000000";
data_b(1205) <= "0000000000";
data_b(1206) <= "0000000000";
data_b(1207) <= "0000000000";
data_b(1208) <= "0000000010";
data_b(1209) <= "0000000010";
data_b(1210) <= "0000000010";
data_b(1211) <= "0000000010";
data_b(1212) <= "0000000000";
data_b(1213) <= "0000000000";
data_b(1214) <= "0000000000";
data_b(1215) <= "0000000000";
-------------------------------------------------------14����
data_b(1216) <= "0000000100";
data_b(1217) <= "0000000100";
data_b(1218) <= "0000000100";
data_b(1219) <= "0000000000";
data_b(1220) <= "0000000000";
data_b(1221) <= "0000000000";
data_b(1222) <= "0000000000";
data_b(1223) <= "0000000000";
data_b(1224) <= "0000000000";
data_b(1225) <= "0000000000";
data_b(1226) <= "0000000000";
data_b(1227) <= "0000000000";
data_b(1228) <= "1000000000";
data_b(1229) <= "1000000000";
data_b(1230) <= "0000000000";
data_b(1231) <= "0000000000";
data_b(1232) <= "0000000000";
data_b(1233) <= "0000000000";
data_b(1234) <= "0000000000";
data_b(1235) <= "0000000000";
data_b(1236) <= "1000000000";
data_b(1237) <= "0000000000";
data_b(1238) <= "0000000000";
data_b(1239) <= "0000000000";
data_b(1240) <= "0000000010";
data_b(1241) <= "0000000010";
data_b(1242) <= "0000000000";
data_b(1243) <= "0000000000";
data_b(1244) <= "0000000000";
data_b(1245) <= "0000000000";
data_b(1246) <= "0000000000";
data_b(1247) <= "0000000000";
------------------------------------------------------15����
data_b(1248) <= "0000000010";                                   
data_b(1249) <= "0000000010";
data_b(1250) <= "0000000010";
data_b(1251) <= "0000000010";
data_b(1252) <= "0000000010";
data_b(1253) <= "0000000010";
data_b(1254) <= "0000000010";
data_b(1255) <= "0000000010";
data_b(1256) <= "0000000010";
data_b(1257) <= "0000000010";
data_b(1258) <= "0000000000";
data_b(1259) <= "0000000000";
data_b(1260) <= "0000000000";
data_b(1261) <= "0000000000";
data_b(1262) <= "0000000000";
data_b(1263) <= "0000000000";
data_b(1264) <= "0000000000";
data_b(1265) <= "0000000000";
data_b(1266) <= "0000000000";
data_b(1267) <= "0000000000";
data_b(1268) <= "1000000000";
data_b(1269) <= "0000000000";
data_b(1270) <= "0000000000";
data_b(1271) <= "0000000000";
data_b(1272) <= "0100000000";
data_b(1273) <= "0000000000";
data_b(1274) <= "0000000000";
data_b(1275) <= "0000000000";
data_b(1276) <= "0010000000";
data_b(1277) <= "0000000000";
data_b(1278) <= "0000000000";
data_b(1279) <= "0000000000";
-------------------------------------------------------16����
data_b(1280) <= "1000000000";          
data_b(1281) <= "1000000000";
data_b(1282) <= "1000000000";
data_b(1283) <= "1000000000";
data_b(1284) <= "1000000000";
data_b(1285) <= "1000000000";
data_b(1286) <= "1000000000";
data_b(1287) <= "1000000000";
data_b(1288) <= "1010000000";
data_b(1289) <= "1000000000";
data_b(1290) <= "1000000000";
data_b(1291) <= "1000000000";
data_b(1292) <= "1000000100";
data_b(1293) <= "1000000000";
data_b(1294) <= "1000000000";
data_b(1295) <= "1000000000";
data_b(1296) <= "0000000010";
data_b(1297) <= "0000000000";
data_b(1298) <= "0000000000";
data_b(1299) <= "0000000000";
data_b(1300) <= "0000000100";
data_b(1301) <= "0000000000";
data_b(1302) <= "0000000000";
data_b(1303) <= "0000000000";
data_b(1304) <= "0000000010";
data_b(1305) <= "0000000000";
data_b(1306) <= "0000000000";
data_b(1307) <= "0000000000";
data_b(1308) <= "0000000001";
data_b(1309) <= "0000000000";
data_b(1310) <= "0000000000";
data_b(1311) <= "0000000000";
---------------------------------------------------------17����
data_b(1312) <= "1000000000";          
data_b(1313) <= "1000000000";
data_b(1314) <= "1000000000";
data_b(1315) <= "1000000000";
data_b(1316) <= "1000000000";
data_b(1317) <= "1000000000";
data_b(1318) <= "1000000000";
data_b(1319) <= "1000000000";
data_b(1320) <= "1010000000";
data_b(1321) <= "1000000000";
data_b(1322) <= "1000000000";
data_b(1323) <= "1000000000";
data_b(1324) <= "1000000100";
data_b(1325) <= "1000000000";
data_b(1326) <= "1000000000";
data_b(1327) <= "1000000000";
data_b(1328) <= "0000000010";
data_b(1329) <= "0000000000";
data_b(1330) <= "0000000000";
data_b(1331) <= "0000000000";
data_b(1332) <= "0000000100";
data_b(1333) <= "0000000000";
data_b(1334) <= "0000000000";
data_b(1335) <= "0000000000";
data_b(1336) <= "0000000010";
data_b(1337) <= "0000000000";
data_b(1338) <= "0000000000";
data_b(1339) <= "0000000000";
data_b(1340) <= "0000000001";
data_b(1341) <= "0000000000";
data_b(1342) <= "0000000000";
data_b(1343) <= "0000000000";
------------------------------------18����
data_b(1344) <= "1000000000";          
data_b(1345) <= "1000000000";
data_b(1346) <= "1000000000";
data_b(1347) <= "1000000000";
data_b(1348) <= "1000000000";
data_b(1349) <= "1000000000";
data_b(1350) <= "1000000000";
data_b(1351) <= "1000000000";
data_b(1352) <= "1010000000";
data_b(1353) <= "1000000000";
data_b(1354) <= "1000000000";
data_b(1355) <= "1000000000";
data_b(1356) <= "1000000100";
data_b(1357) <= "1000000000";
data_b(1358) <= "1000000000";
data_b(1359) <= "1000000000";
data_b(1360) <= "0000000010";
data_b(1361) <= "0000000000";
data_b(1362) <= "0000000000";
data_b(1363) <= "0000000000";
data_b(1364) <= "0000000100";
data_b(1365) <= "0000000000";
data_b(1366) <= "0000000000";
data_b(1367) <= "0000000000";
data_b(1368) <= "0000000010";
data_b(1369) <= "0000000000";
data_b(1370) <= "0000000000";
data_b(1371) <= "0000000000";
data_b(1372) <= "0000000001";
data_b(1373) <= "0000000000";
data_b(1374) <= "0000000000";
data_b(1375) <= "0000000000";
------------------------------------------------------------19����
data_b(1376) <= "1000000000";          
data_b(1377) <= "1000000000";
data_b(1378) <= "1000000000";
data_b(1379) <= "1000000000";
data_b(1380) <= "1000000000";
data_b(1381) <= "1000000000";
data_b(1382) <= "1000000000";
data_b(1383) <= "1000000000";
data_b(1384) <= "1010000000";
data_b(1385) <= "1000000000";
data_b(1386) <= "1000000000";
data_b(1387) <= "1000000000";
data_b(1388) <= "1000000100";
data_b(1389) <= "1000000000";
data_b(1390) <= "1000000000";
data_b(1391) <= "1000000000";
data_b(1392) <= "0000000010";
data_b(1393) <= "0000000000";
data_b(1394) <= "0000000000";
data_b(1395) <= "0000000000";
data_b(1396) <= "0000000100";
data_b(1397) <= "0000000000";
data_b(1398) <= "0000000000";
data_b(1399) <= "0000000000";
data_b(1400) <= "0000000010";
data_b(1401) <= "0000000000";
data_b(1402) <= "0000000000";
data_b(1403) <= "0000000000";
data_b(1404) <= "0000000001";
data_b(1405) <= "0000000000";
data_b(1406) <= "0000000000";
data_b(1407) <= "0000000000";
------------------------------------------------------------------20����
data_b(1408) <= "0000000001";
data_b(1409) <= "0000000000";
data_b(1410) <= "0000000000";
data_b(1411) <= "0000000000";
data_b(1412) <= "0000000001";
data_b(1413) <= "0000000001";
data_b(1414) <= "0000000000";
data_b(1415) <= "0000000000";
data_b(1416) <= "0000000000";
data_b(1417) <= "0000000000";
data_b(1418) <= "0000000000";
data_b(1419) <= "0000000000";
data_b(1420) <= "0000000001";
data_b(1421) <= "0000000001";
data_b(1422) <= "0000000000";
data_b(1423) <= "0000000000";
data_b(1424) <= "0000000000";
data_b(1425) <= "0000000000";
data_b(1426) <= "0000000000";
data_b(1427) <= "0000000000";
data_b(1428) <= "0000000010";
data_b(1429) <= "0000000000";
data_b(1430) <= "0000000000";
data_b(1431) <= "0000000000";
data_b(1432) <= "0000000100";
data_b(1433) <= "0000000100";
data_b(1434) <= "0000000000";
data_b(1435) <= "0000000000";
data_b(1436) <= "0000000000";
data_b(1437) <= "0000000000";
data_b(1438) <= "0000000000";
data_b(1439) <= "0000000000";
------------------------------------21����

data_b(1440) <= "0000000001";
data_b(1441) <= "0000000001";
data_b(1442) <= "0000000001";
data_b(1443) <= "0000000001";
data_b(1444) <= "0000000001";
data_b(1445) <= "0000000001";
data_b(1446) <= "0000000001";
data_b(1447) <= "0000000001";
data_b(1448) <= "0000000001";
data_b(1449) <= "0000000001";
data_b(1450) <= "0000000001";
data_b(1451) <= "0000000001";
data_b(1452) <= "0000000000";
data_b(1453) <= "0000000000";
data_b(1454) <= "0000000000";
data_b(1455) <= "0000000000";
data_b(1456) <= "0000000000";
data_b(1457) <= "0000000000";
data_b(1458) <= "0000000000";
data_b(1459) <= "0000000000";
data_b(1460) <= "0000000000";
data_b(1461) <= "0000000000";
data_b(1462) <= "0000000000";
data_b(1463) <= "0000000000";
data_b(1464) <= "0000000001";
data_b(1465) <= "0000000001";
data_b(1466) <= "0000000000";
data_b(1467) <= "0000000000";
data_b(1468) <= "0000000000";
data_b(1469) <= "0000000000";
data_b(1470) <= "0000000000";
data_b(1471) <= "0000000000";
-----------------------------------------------------------22����
data_b(1472) <= "0000000010";
data_b(1473) <= "0000000010";
data_b(1474) <= "0000000010";
data_b(1475) <= "0000000000";
data_b(1476) <= "0000000000";
data_b(1477) <= "0000000000";
data_b(1478) <= "0000000000";
data_b(1479) <= "0000000000";
data_b(1480) <= "0000000000";
data_b(1481) <= "0000000000";
data_b(1482) <= "0000000000";
data_b(1483) <= "0000000000";
data_b(1484) <= "1000000000";
data_b(1485) <= "1000000000";
data_b(1486) <= "0000000000";
data_b(1487) <= "0000000000";
data_b(1488) <= "0000000000";
data_b(1489) <= "0000000000";
data_b(1490) <= "0000000000";
data_b(1491) <= "0000000000";
data_b(1492) <= "0000000001";
data_b(1493) <= "0000000000";
data_b(1494) <= "0000000000";
data_b(1495) <= "0000000000";
data_b(1496) <= "1000000000";
data_b(1497) <= "0000000000";
data_b(1498) <= "0000000000";
data_b(1499) <= "0000000000";
data_b(1500) <= "0000000001";
data_b(1501) <= "0000000000";
data_b(1502) <= "0000000000";
data_b(1503) <= "0000000000";
-----------------------------------------------------------------23����
data_b(1504) <= "0000000100";
data_b(1505) <= "0000000100";
data_b(1506) <= "0000000100";
data_b(1507) <= "0000000100";
data_b(1508) <= "0000000100";
data_b(1509) <= "0000000100";
data_b(1510) <= "0000000100";
data_b(1511) <= "0000000100";
data_b(1512) <= "0000000100";
data_b(1513) <= "0000000100";
data_b(1514) <= "0000000000";
data_b(1515) <= "0000000000";
data_b(1516) <= "0000000000";
data_b(1517) <= "0000000000";
data_b(1518) <= "0000000000";
data_b(1519) <= "0000000000";
data_b(1520) <= "0000000000";
data_b(1521) <= "0000000000";
data_b(1522) <= "0000000000";
data_b(1523) <= "0000000000";
data_b(1524) <= "1000000000";
data_b(1525) <= "0000000000";
data_b(1526) <= "0000000000";
data_b(1527) <= "0000000000";
data_b(1528) <= "0100000000";
data_b(1529) <= "0000000000";
data_b(1530) <= "0000000000";
data_b(1531) <= "0000000000";
data_b(1532) <= "0010000000";
data_b(1533) <= "0000000000";
data_b(1534) <= "0000000000";
data_b(1535) <= "0000000000";
---------------------------------------24����


----------------------------
--------------------1
scale2(15) <= bm_2;
scale2(16) <= bm_2;
scale2(17) <= bm_2;
scale2(18) <= r;
scale2(19) <= bm_3;
scale2(20) <= bm_3;
scale2(21) <= bm_3;
scale2(22) <= r;
scale2(23) <= bm_2;
scale2(24) <= bm_2;
scale2(25) <= bm_2;
scale2(26) <= r;
scale2(27) <= bm_3;
scale2(28) <= bm_3;
scale2(29) <= bm_3;
scale2(30) <= r;
scale2(31) <= bm_2;
scale2(32) <= bm_2;
scale2(33) <= bm_2;
scale2(34) <= r;
scale2(35) <= bm_3;
scale2(36) <= bm_3;
scale2(37) <= bm_3;
scale2(38) <= r;
scale2(39) <= bm_2;
scale2(40) <= bm_2;
scale2(41) <= bm_2;
scale2(42) <= r;
scale2(43) <= bm_3;
scale2(44) <= bm_3;
scale2(45) <= bm_3;
scale2(46) <= r;
------------------2
scale2(47) <= bm_2;
scale2(48) <= bm_2;
scale2(49) <= bm_2;
scale2(50) <= r;
scale2(51) <= bm_3;
scale2(52) <= bm_3;
scale2(53) <= bm_3;
scale2(54) <= r;
scale2(55) <= bm_2;
scale2(56) <= bm_2;
scale2(57) <= bm_2;
scale2(58) <= r;
scale2(59) <= bm_3;
scale2(60) <= bm_3;
scale2(61) <= bm_3;
scale2(62) <= r;
scale2(63) <= bm_2;
scale2(64) <= bm_2;
scale2(65) <= bm_2;
scale2(66) <= r;
scale2(67) <= bm_3;
scale2(68) <= bm_3;
scale2(69) <= bm_3;
scale2(70) <= r;
scale2(71) <= bm_2;
scale2(72) <= bm_2;
scale2(73) <= bm_2;
scale2(74) <= r;
scale2(75) <= bm_3;
scale2(76) <= bm_3;
scale2(77) <= bm_3;
scale2(78) <= r;
------------------3
scale2(79) <= g_1;
scale2(80) <= g_1;
scale2(81) <= g_1;
scale2(82) <= r;
scale2(83) <= g_2;
scale2(84) <= g_2;
scale2(85) <= g_2;
scale2(86) <= r;
scale2(87) <= g_1;
scale2(88) <= g_1;
scale2(89) <= g_1;
scale2(90) <= r;
scale2(91) <= g_2;
scale2(92) <= g_2;
scale2(93) <= g_2;
scale2(94) <= r;
scale2(95) <= g_1;
scale2(96) <= g_1;
scale2(97) <= g_1;
scale2(98) <= r;
scale2(99) <= g_2;
scale2(100) <= g_2;
scale2(101) <= g_2;
scale2(102) <= r;
scale2(103) <= g_1;
scale2(104) <= g_1;
scale2(105) <= g_1;
scale2(106) <= r;
scale2(107) <= g_2;
scale2(108) <= g_2;
scale2(109) <= g_2;
scale2(110) <= r;
------------------4
scale2(111) <= g_1;
scale2(112) <= g_1;
scale2(113) <= g_1;
scale2(114) <= r;
scale2(115) <= g_2;
scale2(116) <= g_2;
scale2(117) <= g_2;
scale2(118) <= r;
scale2(119) <= g_1;
scale2(120) <= g_1;
scale2(121) <= g_1;
scale2(122) <= r;
scale2(123) <= g_2;
scale2(124) <= g_2;
scale2(125) <= g_2;
scale2(126) <= r;
scale2(127) <= g_1;
scale2(128) <= g_1;
scale2(129) <= g_1;
scale2(130) <= r;
scale2(131) <= g_2;
scale2(132) <= g_2;
scale2(133) <= g_2;
scale2(134) <= r;
scale2(135) <= g_1;
scale2(136) <= g_1;
scale2(137) <= g_1;
scale2(138) <= r;
scale2(139) <= g_2;
scale2(140) <= g_2;
scale2(141) <= g_2;
scale2(142) <= r;
------------------5
scale2(143) <= bm_2;
scale2(144) <= bm_2;
scale2(145) <= bm_2;
scale2(146) <= r;
scale2(147) <= bm_3;
scale2(148) <= bm_3;
scale2(149) <= bm_3;
scale2(150) <= r;
scale2(151) <= bm_2;
scale2(152) <= bm_2;
scale2(153) <= bm_2;
scale2(154) <= r;
scale2(155) <= bm_3;
scale2(156) <= bm_3;
scale2(157) <= bm_3;
scale2(158) <= r;
scale2(159) <= bm_2;
scale2(160) <= bm_2;
scale2(161) <= bm_2;
scale2(162) <= r;
scale2(163) <= bm_3;
scale2(164) <= bm_3;
scale2(165) <= bm_3;
scale2(166) <= r;
scale2(167) <= bm_2;
scale2(168) <= bm_2;
scale2(169) <= bm_2;
scale2(170) <= r;
scale2(171) <= bm_3;
scale2(172) <= bm_3;
scale2(173) <= bm_3;
scale2(174) <= r;
------------------6
scale2(175) <= bm_2;
scale2(176) <= bm_2;
scale2(177) <= bm_2;
scale2(178) <= r;
scale2(179) <= bm_3;
scale2(180) <= bm_3;
scale2(181) <= bm_3;
scale2(182) <= r;
scale2(183) <= bm_2;
scale2(184) <= bm_2;
scale2(185) <= bm_2;
scale2(186) <= r;
scale2(187) <= bm_3;
scale2(188) <= bm_3;
scale2(189) <= bm_3;
scale2(190) <= r;
scale2(191) <= bm_2;
scale2(192) <= bm_2;
scale2(193) <= bm_2;
scale2(194) <= r;
scale2(195) <= bm_3;
scale2(196) <= bm_3;
scale2(197) <= bm_3;
scale2(198) <= r;
scale2(199) <= bm_2;
scale2(200) <= bm_2;
scale2(201) <= bm_2;
scale2(202) <= r;
scale2(203) <= bm_3;
scale2(204) <= bm_3;
scale2(205) <= bm_3;
scale2(206) <= r;
------------------7
scale2(207) <= g_1;
scale2(208) <= g_1;
scale2(209) <= g_1;
scale2(210) <= r;
scale2(211) <= g_2;
scale2(212) <= g_2;
scale2(213) <= g_2;
scale2(214) <= r;
scale2(215) <= g_1;
scale2(216) <= g_1;
scale2(217) <= g_1;
scale2(218) <= r;
scale2(219) <= g_2;
scale2(220) <= g_2;
scale2(221) <= g_2;
scale2(222) <= r;
scale2(223) <= g_1;
scale2(224) <= g_1;
scale2(225) <= g_1;
scale2(226) <= r;
scale2(227) <= g_2;
scale2(228) <= g_2;
scale2(229) <= g_2;
scale2(230) <= r;
scale2(231) <= g_1;
scale2(232) <= g_1;
scale2(233) <= g_1;
scale2(234) <= r;
scale2(235) <= g_2;
scale2(236) <= g_2;
scale2(237) <= g_2;
scale2(238) <= r;
------------------8
scale2(239) <= g_1;
scale2(240) <= g_1;
scale2(241) <= g_1;
scale2(242) <= r;
scale2(243) <= g_2;
scale2(244) <= g_2;
scale2(245) <= g_2;
scale2(246) <= r;
scale2(247) <= g_1;
scale2(248) <= g_1;
scale2(249) <= g_1;
scale2(250) <= r;
scale2(251) <= g_2;
scale2(252) <= g_2;
scale2(253) <= g_2;
scale2(254) <= r;
scale2(255) <= bm_2;
scale2(256) <= bm_2;
scale2(257) <= bm_2;
scale2(258) <= r;
scale2(259) <= f_1;
scale2(260) <= f_1;
scale2(261) <= f_1;
scale2(262) <= r;
scale2(263) <= g_1;
scale2(264) <= g_1;
scale2(265) <= g_1;
scale2(266) <= r;
scale2(267) <= am_1;
scale2(268) <= am_1;
scale2(269) <= am_1;
scale2(270) <= r;
------------------9
scale2(271) <= a_2;
scale2(272) <= a_2;
scale2(273) <= a_2;
scale2(274) <= r;
scale2(275) <= a_3;
scale2(276) <= a_3;
scale2(277) <= a_3;
scale2(278) <= r;
scale2(279) <= a_2;
scale2(280) <= a_2;
scale2(281) <= a_2;
scale2(282) <= r;
scale2(283) <= a_3;
scale2(284) <= a_3;
scale2(285) <= a_3;
scale2(286) <= r;
scale2(287) <= a_2;
scale2(288) <= a_2;
scale2(289) <= a_2;
scale2(290) <= r;
scale2(291) <= f_1;
scale2(292) <= f_1;
scale2(293) <= f_1;
scale2(294) <= r;
scale2(295) <= g_1;
scale2(296) <= g_1;
scale2(297) <= g_1;
scale2(298) <= r;
scale2(299) <= a_2;
scale2(300) <= a_2;
scale2(301) <= a_2;
scale2(302) <= r;
------------------10
scale2(303) <= bm_2;
scale2(304) <= bm_2;
scale2(305) <= bm_2;
scale2(306) <= r;
scale2(307) <= bm_3;
scale2(308) <= bm_3;
scale2(309) <= bm_3;
scale2(310) <= r;
scale2(311) <= bm_2;
scale2(312) <= bm_2;
scale2(313) <= bm_2;
scale2(314) <= r;
scale2(315) <= bm_3;
scale2(316) <= bm_3;
scale2(317) <= bm_3;
scale2(318) <= r;
scale2(319) <= bm_2;
scale2(320) <= bm_2;
scale2(321) <= bm_2;
scale2(322) <= r;
scale2(323) <= f_1;
scale2(324) <= f_1;
scale2(325) <= f_1;
scale2(326) <= r;
scale2(327) <= g_1;
scale2(328) <= g_1;
scale2(329) <= g_1;
scale2(330) <= r;
scale2(331) <= am_1;
scale2(332) <= am_1;
scale2(333) <= am_1;
scale2(334) <= r;
------------------11
scale2(335) <= a_2;
scale2(336) <= a_2;
scale2(337) <= a_2;
scale2(338) <= r;
scale2(339) <= a_3;
scale2(340) <= a_3;
scale2(341) <= a_3;
scale2(342) <= r;
scale2(343) <= a_2;
scale2(344) <= a_2;
scale2(345) <= a_2;
scale2(346) <= r;
scale2(347) <= a_3;
scale2(348) <= a_3;
scale2(349) <= a_3;
scale2(350) <= r;
scale2(351) <= a_2;
scale2(352) <= a_2;
scale2(353) <= a_2;
scale2(354) <= r;
scale2(355) <= f_1;
scale2(356) <= f_1;
scale2(357) <= f_1;
scale2(358) <= r;
scale2(359) <= g_1;
scale2(360) <= g_1;
scale2(361) <= g_1;
scale2(362) <= r;
scale2(363) <= a_2;
scale2(364) <= a_2;
scale2(365) <= a_2;
scale2(366) <= r;
-------------------12
scale2(367) <= bm_2;
scale2(368) <= bm_2;
scale2(369) <= bm_2;
scale2(370) <= r;
scale2(371) <= bm_3;
scale2(372) <= bm_3;
scale2(373) <= bm_3;
scale2(374) <= r;
scale2(375) <= bm_2;
scale2(376) <= bm_2;
scale2(377) <= bm_2;
scale2(378) <= r;
scale2(379) <= bm_3;
scale2(380) <= bm_3;
scale2(381) <= bm_3;
scale2(382) <= r;
scale2(383) <= bm_2;
scale2(384) <= bm_2;
scale2(385) <= bm_2;
scale2(386) <= r;
scale2(387) <= bm_2;
scale2(388) <= bm_2;
scale2(389) <= bm_2;
scale2(390) <= r;
scale2(391) <= c_2;
scale2(392) <= c_2;
scale2(393) <= c_2;
scale2(394) <= r;
scale2(395) <= d_2;
scale2(396) <= d_2;
scale2(397) <= d_2;
scale2(398) <= r;
------------------13
scale2(399) <= em_2;
scale2(400) <= em_2;
scale2(401) <= em_2;
scale2(402) <= r;
scale2(403) <= em_3;
scale2(404) <= em_3;
scale2(405) <= em_3;
scale2(406) <= r;
scale2(407) <= em_2;
scale2(408) <= em_2;
scale2(409) <= em_2;
scale2(410) <= r;
scale2(411) <= em_3;
scale2(412) <= em_3;
scale2(413) <= em_3;
scale2(414) <= r;
scale2(415) <= em_2;
scale2(416) <= em_2;
scale2(417) <= em_2;
scale2(418) <= r;
scale2(419) <= em_3;
scale2(420) <= em_3;
scale2(421) <= em_3;
scale2(422) <= r;
scale2(423) <= em_2;
scale2(424) <= em_2;
scale2(425) <= em_2;
scale2(426) <= r;
scale2(427) <= em_3;
scale2(428) <= em_3;
scale2(429) <= em_3;
scale2(430) <= r;
------------------14
scale2(431) <= d_2;
scale2(432) <= d_2;
scale2(433) <= d_2;
scale2(434) <= r;
scale2(435) <= d_3;
scale2(436) <= d_3;
scale2(437) <= d_3;
scale2(438) <= r;
scale2(439) <= d_2;
scale2(440) <= d_2;
scale2(441) <= d_2;
scale2(442) <= r;
scale2(443) <= d_3;
scale2(444) <= d_3;
scale2(445) <= d_3;
scale2(446) <= r;
scale2(447) <= d_2;
scale2(448) <= d_2;
scale2(449) <= d_2;
scale2(450) <= r;
scale2(451) <= d_3;
scale2(452) <= d_3;
scale2(453) <= d_3;
scale2(454) <= r;
scale2(455) <= d_2;
scale2(456) <= d_2;
scale2(457) <= d_2;
scale2(458) <= r;
scale2(459) <= d_3;
scale2(460) <= d_3;
scale2(461) <= d_3;
scale2(462) <= r;
------------------15
scale2(463) <= c_2;
scale2(464) <= c_2;
scale2(465) <= c_2;
scale2(466) <= r;
scale2(467) <= c_3;
scale2(468) <= c_3;
scale2(469) <= c_3;
scale2(470) <= r;
scale2(471) <= c_2;
scale2(472) <= c_2;
scale2(473) <= c_2;
scale2(474) <= r;
scale2(475) <= c_3;
scale2(476) <= c_3;
scale2(477) <= c_3;
scale2(478) <= r;
scale2(479) <= g_1;
scale2(480) <= g_1;
scale2(481) <= g_1;
scale2(482) <= r;
scale2(483) <= g_2;
scale2(484) <= g_2;
scale2(485) <= g_2;
scale2(486) <= r;
scale2(487) <= g_1;
scale2(488) <= g_1;
scale2(489) <= g_1;
scale2(490) <= r;
scale2(491) <= g_2;
scale2(492) <= g_2;
scale2(493) <= g_2;
scale2(494) <= r;
------------------16
scale2(495) <= c_2;
scale2(496) <= c_2;
scale2(497) <= c_2;
scale2(498) <= r;
scale2(499) <= c_3;
scale2(500) <= c_3;
scale2(501) <= c_3;
scale2(502) <= r;
scale2(503) <= c_2;
scale2(504) <= c_2;
scale2(505) <= c_2;
scale2(506) <= r;
scale2(507) <= c_3;
scale2(508) <= c_3;
scale2(509) <= c_3;
scale2(510) <= r;
scale2(511) <= c_2;
scale2(512) <= c_2;
scale2(513) <= c_2;
scale2(514) <= r;
scale2(515) <= f_1;
scale2(516) <= f_1;
scale2(517) <= f_1;
scale2(518) <= r;
scale2(519) <= g_1;
scale2(520) <= g_1;
scale2(521) <= g_1;
scale2(522) <= r;
scale2(523) <= am_1;
scale2(524) <= am_1;
scale2(525) <= am_1; 
scale2(526) <= r;
------------------17
scale2(527) <= a_2;
scale2(528) <= a_2;
scale2(529) <= a_2;
scale2(530) <= r;
scale2(531) <= a_3;
scale2(532) <= a_3;
scale2(533) <= a_3;
scale2(534) <= r;
scale2(535) <= a_2;
scale2(536) <= a_2;
scale2(537) <= a_2;
scale2(538) <= r;
scale2(539) <= a_3;
scale2(540) <= a_3;
scale2(541) <= a_3;
scale2(542) <= r;
scale2(543) <= a_2;
scale2(544) <= a_2;
scale2(545) <= a_2;
scale2(546) <= r;
scale2(547) <= f_1;
scale2(548) <= f_1;
scale2(549) <= f_1;
scale2(550) <= r;
scale2(551) <= g_1;
scale2(552) <= g_1;
scale2(553) <= g_1;
scale2(554) <= r;
scale2(555) <= a_2;
scale2(556) <= a_2;
scale2(557) <= a_2;
scale2(558) <= r;
------------------18
scale2(559) <= bm_2;
scale2(560) <= bm_2;
scale2(561) <= bm_2;
scale2(562) <= r;
scale2(563) <= bm_3;
scale2(564) <= bm_3;
scale2(565) <= bm_3;
scale2(566) <= r;
scale2(567) <= bm_2;
scale2(568) <= bm_2;
scale2(569) <= bm_2;
scale2(570) <= r;
scale2(571) <= bm_3;
scale2(572) <= bm_3;
scale2(573) <= bm_3;
scale2(574) <= r;
scale2(575) <= bm_2;
scale2(576) <= bm_2;
scale2(577) <= bm_2;
scale2(578) <= r;
scale2(579) <= f_1;
scale2(580) <= f_1;
scale2(581) <= f_1;
scale2(582) <= r;
scale2(583) <= g_1;
scale2(584) <= g_1;
scale2(585) <= g_1;
scale2(586) <= r;
scale2(587) <= am_1;
scale2(588) <= am_1;
scale2(589) <= am_1;
scale2(590) <= r;
------------------19
scale2(591) <= a_2;
scale2(592) <= a_2;
scale2(593) <= a_2;
scale2(594) <= r;
scale2(595) <= a_3;
scale2(596) <= a_3;
scale2(597) <= a_3;
scale2(598) <= r;
scale2(599) <= a_2;
scale2(600) <= a_2;
scale2(601) <= a_2;
scale2(602) <= r;
scale2(603) <= a_3;
scale2(604) <= a_3;
scale2(605) <= a_3;
scale2(606) <= r;
scale2(607) <= a_2;
scale2(608) <= a_2;
scale2(609) <= a_2;
scale2(610) <= r;
scale2(611) <= f_1;
scale2(612) <= f_1;
scale2(613) <= f_1;
scale2(614) <= r;
scale2(615) <= g_1;
scale2(616) <= g_1;
scale2(617) <= g_1;
scale2(618) <= r;
scale2(619) <= a_2;
scale2(620) <= a_2;
scale2(621) <= a_2;
scale2(622) <= r;
-------------------20
scale2(623) <= bm_2;
scale2(624) <= bm_2;
scale2(625) <= bm_2;
scale2(626) <= r;
scale2(627) <= bm_3;
scale2(628) <= bm_3;
scale2(629) <= bm_3;
scale2(630) <= r;
scale2(631) <= bm_2;
scale2(632) <= bm_2;
scale2(633) <= bm_2;
scale2(634) <= r;
scale2(635) <= bm_3;
scale2(636) <= bm_3;
scale2(637) <= bm_3;
scale2(638) <= r;
scale2(639) <= bm_2;
scale2(640) <= bm_2;
scale2(641) <= bm_2;
scale2(642) <= r;
scale2(643) <= bm_2;
scale2(644) <= bm_2;
scale2(645) <= bm_2;
scale2(646) <= r;
scale2(647) <= c_2;
scale2(648) <= c_2;
scale2(649) <= c_2;
scale2(650) <= r;
scale2(651) <= d_2;
scale2(652) <= d_2;
scale2(653) <= d_2;
scale2(654) <= r;
------------------21
scale2(655) <= em_2;
scale2(656) <= em_2;
scale2(657) <= em_2;
scale2(658) <= r;
scale2(659) <= em_3;
scale2(660) <= em_3;
scale2(661) <= em_3;
scale2(662) <= r;
scale2(663) <= em_2;
scale2(664) <= em_2;
scale2(665) <= em_2;
scale2(666) <= r;
scale2(667) <= em_3;
scale2(668) <= em_3;
scale2(669) <= em_3;
scale2(670) <= r;
scale2(671) <= em_2;
scale2(672) <= em_2;
scale2(673) <= em_2;
scale2(674) <= r;
scale2(675) <= em_3;
scale2(676) <= em_3;
scale2(677) <= em_3;
scale2(678) <= r;
scale2(679) <= em_2;
scale2(680) <= em_2;
scale2(681) <= em_2;
scale2(682) <= r;
scale2(683) <= em_3;
scale2(684) <= em_3;
scale2(685) <= em_3;
scale2(686) <= r;
------------------22
scale2(687) <= d_2;
scale2(688) <= d_2;
scale2(689) <= d_2;
scale2(690) <= r;
scale2(691) <= d_3;
scale2(692) <= d_3;
scale2(693) <= d_3;
scale2(694) <= r;
scale2(695) <= d_2;
scale2(696) <= d_2;
scale2(697) <= d_2;
scale2(698) <= r;
scale2(699) <= d_3;
scale2(700) <= d_3;
scale2(701) <= d_3;
scale2(702) <= r;
scale2(703) <= d_2;
scale2(704) <= d_2;
scale2(705) <= d_2;
scale2(706) <= r;
scale2(707) <= d_3;
scale2(708) <= d_3;
scale2(709) <= d_3;
scale2(710) <= r;
scale2(711) <= d_2;
scale2(712) <= d_2;
scale2(713) <= d_2;
scale2(714) <= r;
scale2(715) <= d_3;
scale2(716) <= d_3;
scale2(717) <= d_3;
scale2(718) <= r;
------------------23
scale2(719) <= c_2;
scale2(720) <= c_2;
scale2(721) <= c_2;
scale2(722) <= r;
scale2(723) <= c_3;
scale2(724) <= c_3;
scale2(725) <= c_3;
scale2(726) <= r;
scale2(727) <= c_2;
scale2(728) <= c_2;
scale2(729) <= c_2;
scale2(730) <= r;
scale2(731) <= c_3;
scale2(732) <= c_3;
scale2(733) <= c_3;
scale2(734) <= r;
scale2(735) <= f_1;
scale2(736) <= f_1;
scale2(737) <= f_1;
scale2(738) <= r;
scale2(739) <= c_2;
scale2(740) <= c_2;
scale2(741) <= c_2;
scale2(742) <= r;
scale2(743) <= f_1;
scale2(744) <= f_1;
scale2(745) <= f_1;
scale2(746) <= r;
scale2(747) <= c_2;
scale2(748) <= c_2;
scale2(749) <= c_2;
scale2(750) <= r;
------------------24
scale2(751) <= bm_2;
scale2(752) <= bm_2;
scale2(753) <= bm_2;
scale2(754) <= bm_2;
scale2(755) <= bm_2;
scale2(756) <= bm_2;
scale2(757) <= bm_2;
scale2(758) <= bm_2;
scale2(759) <= bm_2;
scale2(760) <= bm_2;
scale2(761) <= bm_2;
scale2(762) <= bm_2;
scale2(763) <= bm_2;
scale2(764) <= bm_2;
scale2(765) <= bm_2;
scale2(766) <= bm_2;
scale2(767) <= bm_2;
scale2(768) <= bm_2;
scale2(769) <= bm_2;
scale2(770) <= r;
scale2(771) <= f_1;
scale2(772) <= f_1;
scale2(773) <= f_1;
scale2(774) <= r;
scale2(775) <= g_1;
scale2(776) <= g_1;
scale2(777) <= g_1;
scale2(778) <= r;
scale2(779) <= a_2;
scale2(780) <= a_2;
scale2(781) <= a_2;
scale2(782) <= r;
------------------25
scale2(783) <= bm_2;
scale2(784) <= bm_2;
scale2(785) <= bm_2;
scale2(786) <= r;
scale2(787) <= bm_3;
scale2(788) <= bm_3;
scale2(789) <= bm_3;
scale2(790) <= r;
scale2(791) <= bm_2;
scale2(792) <= bm_2;
scale2(793) <= bm_2;
scale2(794) <= r;
scale2(795) <= bm_3;
scale2(796) <= bm_3;
scale2(797) <= bm_3;
scale2(798) <= r;
scale2(799) <= bm_2;
scale2(800) <= bm_2;
scale2(801) <= bm_2;
scale2(802) <= r;
scale2(803) <= bm_3;
scale2(804) <= bm_3;
scale2(805) <= bm_3;
scale2(806) <= r;
scale2(807) <= bm_2;
scale2(808) <= bm_2;
scale2(809) <= bm_2;
scale2(810) <= r;
scale2(811) <= bm_3;
scale2(812) <= bm_3;
scale2(813) <= bm_3;
scale2(814) <= r;
------------------26
scale2(815) <= bm_2;
scale2(816) <= bm_2;
scale2(817) <= bm_2;
scale2(818) <= r;
scale2(819) <= bm_3;
scale2(820) <= bm_3;
scale2(821) <= bm_3;
scale2(822) <= r;
scale2(823) <= bm_2;
scale2(824) <= bm_2;
scale2(825) <= bm_2;
scale2(826) <= r;
scale2(827) <= bm_3;
scale2(828) <= bm_3;
scale2(829) <= bm_3;
scale2(830) <= r;
scale2(831) <= bm_2;
scale2(832) <= bm_2;
scale2(833) <= bm_2;
scale2(834) <= r;
scale2(835) <= bm_3;
scale2(836) <= bm_3;
scale2(837) <= bm_3;
scale2(838) <= r;
scale2(839) <= bm_2;
scale2(840) <= bm_2;
scale2(841) <= bm_2;
scale2(842) <= r;
scale2(843) <= bm_3;
scale2(844) <= bm_3;
scale2(845) <= bm_3;
scale2(846) <= r;
------------------27
scale2(847) <= g_1;
scale2(848) <= g_1;
scale2(849) <= g_1;
scale2(850) <= r;
scale2(851) <= g_2;
scale2(852) <= g_2;
scale2(853) <= g_2;
scale2(854) <= r;
scale2(855) <= g_1;
scale2(856) <= g_1;
scale2(857) <= g_1;
scale2(858) <= r;
scale2(859) <= g_2;
scale2(860) <= g_2;
scale2(861) <= g_2;
scale2(862) <= r;
scale2(863) <= g_1;
scale2(864) <= g_1;
scale2(865) <= g_1;
scale2(866) <= r;
scale2(867) <= g_2;
scale2(868) <= g_2;
scale2(869) <= g_2;
scale2(870) <= r;
scale2(871) <= g_1;
scale2(872) <= g_1;
scale2(873) <= g_1;
scale2(874) <= r;
scale2(875) <= g_2;
scale2(876) <= g_2;
scale2(877) <= g_2;
scale2(878) <= r;
------------------28
scale2(879) <= g_1;
scale2(880) <= g_1;
scale2(881) <= g_1;
scale2(882) <= r;
scale2(883) <= g_2;
scale2(884) <= g_2;
scale2(885) <= g_2;
scale2(886) <= r;
scale2(887) <= g_1;
scale2(888) <= g_1;
scale2(889) <= g_1;
scale2(890) <= r;
scale2(891) <= g_2;
scale2(892) <= g_2;
scale2(893) <= g_2;
scale2(894) <= r;
scale2(895) <= g_1;
scale2(896) <= g_1;
scale2(897) <= g_1;
scale2(898) <= r;
scale2(899) <= g_2;
scale2(900) <= g_2;
scale2(901) <= g_2;
scale2(902) <= r;
scale2(903) <= g_1;
scale2(904) <= g_1;
scale2(905) <= g_1;
scale2(906) <= r;
scale2(907) <= g_2;
scale2(908) <= g_2;
scale2(909) <= g_2;
scale2(910) <= r;
------------------29
scale2(911) <= bm_2;
scale2(912) <= bm_2;
scale2(913) <= bm_2;
scale2(914) <= r;
scale2(915) <= bm_3;
scale2(916) <= bm_3;
scale2(917) <= bm_3;
scale2(918) <= r;
scale2(919) <= bm_2;
scale2(920) <= bm_2;
scale2(921) <= bm_2;
scale2(922) <= r;
scale2(923) <= bm_3;
scale2(924) <= bm_3;
scale2(925) <= bm_3;
scale2(926) <= r;
scale2(927) <= bm_2;
scale2(928) <= bm_2;
scale2(929) <= bm_2;
scale2(930) <= r;
scale2(931) <= bm_3;
scale2(932) <= bm_3;
scale2(933) <= bm_3;
scale2(934) <= r;
scale2(935) <= bm_2;
scale2(936) <= bm_2;
scale2(937) <= bm_2;
scale2(938) <= r;
scale2(939) <= bm_3;
scale2(940) <= bm_3;
scale2(941) <= bm_3;
scale2(942) <= r;
------------------30
scale2(943) <= bm_2;
scale2(944) <= bm_2;
scale2(945) <= bm_2;
scale2(946) <= r;
scale2(947) <= bm_3;
scale2(948) <= bm_3;
scale2(949) <= bm_3;
scale2(950) <= r;
scale2(951) <= bm_2;
scale2(952) <= bm_2;
scale2(953) <= bm_2;
scale2(954) <= r;
scale2(955) <= bm_3;
scale2(956) <= bm_3;
scale2(957) <= bm_3;
scale2(958) <= r;
scale2(959) <= bm_2;
scale2(960) <= bm_2;
scale2(961) <= bm_2;
scale2(962) <= r;
scale2(963) <= bm_3;
scale2(964) <= bm_3;
scale2(965) <= bm_3;
scale2(966) <= r;
scale2(967) <= bm_2;
scale2(968) <= bm_2;
scale2(969) <= bm_2;
scale2(970) <= r;
scale2(971) <= bm_3;
scale2(972) <= bm_3;
scale2(973) <= bm_3;
scale2(974) <= r;
------------------31
scale2(975) <= g_1;
scale2(976) <= g_1;
scale2(977) <= g_1;
scale2(978) <= r;
scale2(979) <= g_2;
scale2(980) <= g_2;
scale2(981) <= g_2;
scale2(982) <= r;
scale2(983) <= g_1;
scale2(984) <= g_1;
scale2(985) <= g_1;
scale2(986) <= r;
scale2(987) <= g_2;
scale2(988) <= g_2;
scale2(989) <= g_2;
scale2(990) <= r;
scale2(991) <= g_1;
scale2(992) <= g_1;
scale2(993) <= g_1;
scale2(994) <= r;
scale2(995) <= g_2;
scale2(996) <= g_2;
scale2(997) <= g_2;
scale2(998) <= r;
scale2(999) <= g_1;
scale2(1000) <= g_1;
scale2(1001) <= g_1;
scale2(1002) <= r;
scale2(1003) <= g_2;
scale2(1004) <= g_2;
scale2(1005) <= g_2;
scale2(1006) <= r;
------------------32
scale2(1007) <= g_1;
scale2(1008) <= g_1;
scale2(1009) <= g_1;
scale2(1010) <= r;
scale2(1011) <= g_2;
scale2(1012) <= g_2;
scale2(1013) <= g_2;
scale2(1014) <= r;
scale2(1015) <= g_1;
scale2(1016) <= g_1;
scale2(1017) <= g_1;
scale2(1018) <= r;
scale2(1019) <= g_2;
scale2(1020) <= g_2;
scale2(1021) <= g_2;
scale2(1022) <= r;
scale2(1023) <= bm_2;
scale2(1024) <= bm_2;
scale2(1025) <= bm_2;
scale2(1026) <= r;
scale2(1027) <= f_1;
scale2(1028) <= f_1;
scale2(1029) <= f_1;
scale2(1030) <= r;
scale2(1031) <= g_1;
scale2(1032) <= g_1;
scale2(1033) <= g_1;
scale2(1034) <= r;
scale2(1035) <= am_1;
scale2(1036) <= am_1;
scale2(1037) <= am_1;
scale2(1038) <= r;
------------------33
scale2(1039) <= a_2;
scale2(1040) <= a_2;
scale2(1041) <= a_2;
scale2(1042) <= r;
scale2(1043) <= a_3;
scale2(1044) <= a_3;
scale2(1045) <= a_3;
scale2(1046) <= r;
scale2(1047) <= a_2;
scale2(1048) <= a_2;
scale2(1049) <= a_2;
scale2(1050) <= r;
scale2(1051) <= a_3;
scale2(1052) <= a_3;
scale2(1053) <= a_3;
scale2(1054) <= r;
scale2(1055) <= a_2;
scale2(1056) <= a_2;
scale2(1057) <= a_2;
scale2(1058) <= r;
scale2(1059) <= f_1;
scale2(1060) <= f_1;
scale2(1061) <= f_1;
scale2(1062) <= r;
scale2(1063) <= g_1;
scale2(1064) <= g_1;
scale2(1065) <= g_1;
scale2(1066) <= r;
scale2(1067) <= a_2;
scale2(1068) <= a_2;
scale2(1069) <= a_2;
scale2(1070) <= r;
------------------34
scale2(1071) <= bm_2;
scale2(1072) <= bm_2;
scale2(1073) <= bm_2;
scale2(1074) <= r;
scale2(1075) <= bm_3;
scale2(1076) <= bm_3;
scale2(1077) <= bm_3;
scale2(1078) <= r;
scale2(1079) <= bm_2;
scale2(1080) <= bm_2;
scale2(1081) <= bm_2;
scale2(1082) <= r;
scale2(1083) <= bm_3;
scale2(1084) <= bm_3;
scale2(1085) <= bm_3;
scale2(1086) <= r;
scale2(1087) <= bm_2;
scale2(1088) <= bm_2;
scale2(1089) <= bm_2;
scale2(1090) <= r;
scale2(1091) <= f_1;
scale2(1092) <= f_1;
scale2(1093) <= f_1;
scale2(1094) <= r;
scale2(1095) <= g_1;
scale2(1096) <= g_1;
scale2(1097) <= g_1;
scale2(1098) <= r;
scale2(1099) <= am_1;
scale2(1100) <= am_1;
scale2(1101) <= am_1;
scale2(1102) <= r;
------------------35
scale2(1103) <= a_2;
scale2(1104) <= a_2;
scale2(1105) <= a_2;
scale2(1106) <= r;
scale2(1107) <= a_3;
scale2(1108) <= a_3;
scale2(1109) <= a_3;
scale2(1110) <= r;
scale2(1111) <= a_2;
scale2(1112) <= a_2;
scale2(1113) <= a_2;
scale2(1114) <= r;
scale2(1115) <= a_3;
scale2(1116) <= a_3;
scale2(1117) <= a_3;
scale2(1118) <= r;
scale2(1119) <= a_2;
scale2(1120) <= a_2;
scale2(1121) <= a_2;
scale2(1122) <= r;
scale2(1123) <= f_1;
scale2(1124) <= f_1;
scale2(1125) <= f_1;
scale2(1126) <= r;
scale2(1127) <= g_1;
scale2(1128) <= g_1;
scale2(1129) <= g_1;
scale2(1130) <= r;
scale2(1131) <= a_2;
scale2(1132) <= a_2;
scale2(1133) <= a_2;
scale2(1134) <= r;
-------------------36
scale2(1135) <= bm_2;
scale2(1136) <= bm_2;
scale2(1137) <= bm_2;
scale2(1138) <= r;
scale2(1139) <= bm_3;
scale2(1140) <= bm_3;
scale2(1141) <= bm_3;
scale2(1142) <= r;
scale2(1143) <= bm_2;
scale2(1144) <= bm_2;
scale2(1145) <= bm_2;
scale2(1146) <= r;
scale2(1147) <= bm_3;
scale2(1148) <= bm_3;
scale2(1149) <= bm_3;
scale2(1150) <= r;
scale2(1151) <= bm_2;
scale2(1152) <= bm_2;
scale2(1153) <= bm_2;
scale2(1154) <= r;
scale2(1155) <= bm_2;
scale2(1156) <= bm_2;
scale2(1157) <= bm_2;
scale2(1158) <= r;
scale2(1159) <= c_2;
scale2(1160) <= c_2;
scale2(1161) <= c_2;
scale2(1162) <= r;
scale2(1163) <= d_2;
scale2(1164) <= d_2;
scale2(1165) <= d_2;
scale2(1166) <= r;
------------------37
scale2(1167) <= em_2;
scale2(1168) <= em_2;
scale2(1169) <= em_2;
scale2(1170) <= r;
scale2(1171) <= em_3;
scale2(1172) <= em_3;
scale2(1173) <= em_3;
scale2(1174) <= r;
scale2(1175) <= em_2;
scale2(1176) <= em_2;
scale2(1177) <= em_2;
scale2(1178) <= r;
scale2(1179) <= em_3;
scale2(1180) <= em_3;
scale2(1181) <= em_3;
scale2(1182) <= r;
scale2(1183) <= em_2;
scale2(1184) <= em_2;
scale2(1185) <= em_2;
scale2(1186) <= r;
scale2(1187) <= em_3;
scale2(1188) <= em_3;
scale2(1189) <= em_3;
scale2(1190) <= r;
scale2(1191) <= em_2;
scale2(1192) <= em_2;
scale2(1193) <= em_2;
scale2(1194) <= r;
scale2(1195) <= em_3;
scale2(1196) <= em_3;
scale2(1197) <= em_3;
scale2(1198) <= r;
------------------38
scale2(1199) <= d_2;
scale2(1200) <= d_2;
scale2(1201) <= d_2;
scale2(1202) <= r;
scale2(1203) <= d_3;
scale2(1204) <= d_3;
scale2(1205) <= d_3;
scale2(1206) <= r;
scale2(1207) <= d_2;
scale2(1208) <= d_2;
scale2(1209) <= d_2;
scale2(1210) <= r;
scale2(1211) <= d_3;
scale2(1212) <= d_3;
scale2(1213) <= d_3;
scale2(1214) <= r;
scale2(1215) <= d_2;
scale2(1216) <= d_2;
scale2(1217) <= d_2;
scale2(1218) <= r;
scale2(1219) <= d_3;
scale2(1220) <= d_3;
scale2(1221) <= d_3;
scale2(1222) <= r;
scale2(1223) <= d_2;
scale2(1224) <= d_2;
scale2(1225) <= d_2;
scale2(1226) <= r;
scale2(1227) <= d_3;
scale2(1228) <= d_3;
scale2(1229) <= d_3;
scale2(1230) <= r;
------------------39
scale2(1231) <= c_2;
scale2(1232) <= c_2;
scale2(1233) <= c_2;
scale2(1234) <= r;
scale2(1235) <= c_3;
scale2(1236) <= c_3;
scale2(1237) <= c_3;
scale2(1238) <= r;
scale2(1239) <= c_2;
scale2(1240) <= c_2;
scale2(1241) <= c_2;
scale2(1242) <= r;
scale2(1243) <= c_3;
scale2(1244) <= c_3;
scale2(1245) <= c_3;
scale2(1246) <= r;
scale2(1247) <= g_1;
scale2(1248) <= g_1;
scale2(1249) <= g_1;
scale2(1250) <= r;
scale2(1251) <= g_2;
scale2(1252) <= g_2;
scale2(1253) <= g_2;
scale2(1254) <= r;
scale2(1255) <= g_1;
scale2(1256) <= g_1;
scale2(1257) <= g_1;
scale2(1258) <= r;
scale2(1259) <= g_2;
scale2(1260) <= g_2;
scale2(1261) <= g_2;
scale2(1262) <= r;
------------------40
scale2(1263) <= c_2;
scale2(1264) <= c_2;
scale2(1265) <= c_2;
scale2(1266) <= r;
scale2(1267) <= c_3;
scale2(1268) <= c_3;
scale2(1269) <= c_3;
scale2(1270) <= r;
scale2(1271) <= c_2;
scale2(1272) <= c_2;
scale2(1273) <= c_2;
scale2(1274) <= r;
scale2(1275) <= c_3;
scale2(1276) <= c_3;
scale2(1277) <= c_3;
scale2(1278) <= r;
scale2(1279) <= c_2;
scale2(1280) <= c_2;
scale2(1281) <= c_2;
scale2(1282) <= r;
scale2(1283) <= f_1;
scale2(1284) <= f_1;
scale2(1285) <= f_1;
scale2(1286) <= r;
scale2(1287) <= g_1;
scale2(1288) <= g_1;
scale2(1289) <= g_1;
scale2(1290) <= r;
scale2(1291) <= am_1;
scale2(1292) <= am_1;
scale2(1293) <= am_1; 
scale2(1294) <= r;
------------------41
scale2(1295) <= a_2;
scale2(1296) <= a_2;
scale2(1297) <= a_2;
scale2(1298) <= r;
scale2(1299) <= a_3;
scale2(1300) <= a_3;
scale2(1301) <= a_3;
scale2(1302) <= r;
scale2(1303) <= a_2;
scale2(1304) <= a_2;
scale2(1305) <= a_2;
scale2(1306) <= r;
scale2(1307) <= a_3;
scale2(1308) <= a_3;
scale2(1309) <= a_3;
scale2(1310) <= r;
scale2(1311) <= a_2;
scale2(1312) <= a_2;
scale2(1313) <= a_2;
scale2(1314) <= r;
scale2(1315) <= f_1;
scale2(1316) <= f_1;
scale2(1317) <= f_1;
scale2(1318) <= r;
scale2(1319) <= g_1;
scale2(1320) <= g_1;
scale2(1321) <= g_1;
scale2(1322) <= r;
scale2(1323) <= a_2;
scale2(1324) <= a_2;
scale2(1325) <= a_2;
scale2(1326) <= r;
------------------42
scale2(1327) <= bm_2;
scale2(1328) <= bm_2;
scale2(1329) <= bm_2;
scale2(1330) <= r;
scale2(1331) <= bm_3;
scale2(1332) <= bm_3;
scale2(1333) <= bm_3;
scale2(1334) <= r;
scale2(1335) <= bm_2;
scale2(1336) <= bm_2;
scale2(1337) <= bm_2;
scale2(1338) <= r;
scale2(1339) <= bm_3;
scale2(1340) <= bm_3;
scale2(1341) <= bm_3;
scale2(1342) <= r;
scale2(1343) <= bm_2;
scale2(1344) <= bm_2;
scale2(1345) <= bm_2;
scale2(1346) <= r;
scale2(1347) <= f_1;
scale2(1348) <= f_1;
scale2(1349) <= f_1;
scale2(1350) <= r;
scale2(1351) <= g_1;
scale2(1352) <= g_1;
scale2(1353) <= g_1;
scale2(1354) <= r;
scale2(1355) <= am_1;
scale2(1356) <= am_1;
scale2(1357) <= am_1;
scale2(1358) <= r;
------------------43
scale2(1359) <= a_2;
scale2(1360) <= a_2;
scale2(1361) <= a_2;
scale2(1362) <= r;
scale2(1363) <= a_3;
scale2(1364) <= a_3;
scale2(1365) <= a_3;
scale2(1366) <= r;
scale2(1367) <= a_2;
scale2(1368) <= a_2;
scale2(1369) <= a_2;
scale2(1370) <= r;
scale2(1371) <= a_3;
scale2(1372) <= a_3;
scale2(1373) <= a_3;
scale2(1374) <= r;
scale2(1375) <= a_2;
scale2(1376) <= a_2;
scale2(1377) <= a_2;
scale2(1378) <= r;
scale2(1379) <= f_1;
scale2(1380) <= f_1;
scale2(1381) <= f_1;
scale2(1382) <= r;
scale2(1383) <= g_1;
scale2(1384) <= g_1;
scale2(1385) <= g_1;
scale2(1386) <= r;
scale2(1387) <= a_2;
scale2(1388) <= a_2;
scale2(1389) <= a_2;
scale2(1390) <= r;
-------------------44
scale2(1391) <= bm_2;
scale2(1392) <= bm_2;
scale2(1393) <= bm_2;
scale2(1394) <= r;
scale2(1395) <= bm_3;
scale2(1396) <= bm_3;
scale2(1397) <= bm_3;
scale2(1398) <= r;
scale2(1399) <= bm_2;
scale2(1400) <= bm_2;
scale2(1401) <= bm_2;
scale2(1402) <= r;
scale2(1403) <= bm_3;
scale2(1404) <= bm_3;
scale2(1405) <= bm_3;
scale2(1406) <= r;
scale2(1407) <= bm_2;
scale2(1408) <= bm_2;
scale2(1409) <= bm_2;
scale2(1410) <= r;
scale2(1411) <= bm_2;
scale2(1412) <= bm_2;
scale2(1413) <= bm_2;
scale2(1414) <= r;
scale2(1415) <= c_2;
scale2(1416) <= c_2;
scale2(1417) <= c_2;
scale2(1418) <= r;
scale2(1419) <= d_2;
scale2(1420) <= d_2;
scale2(1421) <= d_2;
scale2(1422) <= r;
------------------45
scale2(1423) <= em_2;
scale2(1424) <= em_2;
scale2(1425) <= em_2;
scale2(1426) <= r;
scale2(1427) <= em_3;
scale2(1428) <= em_3;
scale2(1429) <= em_3;
scale2(1430) <= r;
scale2(1431) <= em_2;
scale2(1432) <= em_2;
scale2(1433) <= em_2;
scale2(1434) <= r;
scale2(1435) <= em_3;
scale2(1436) <= em_3;
scale2(1437) <= em_3;
scale2(1438) <= r;
scale2(1439) <= em_2;
scale2(1440) <= em_2;
scale2(1441) <= em_2;
scale2(1442) <= r;
scale2(1443) <= em_3;
scale2(1444) <= em_3;
scale2(1445) <= em_3;
scale2(1446) <= r;
scale2(1447) <= em_2;
scale2(1448) <= em_2;
scale2(1449) <= em_2;
scale2(1450) <= r;
scale2(1451) <= em_3;
scale2(1452) <= em_3;
scale2(1453) <= em_3;
scale2(1454) <= r;
------------------46
scale2(1455) <= d_2;
scale2(1456) <= d_2;
scale2(1457) <= d_2;
scale2(1458) <= r;
scale2(1459) <= d_3;
scale2(1460) <= d_3;
scale2(1461) <= d_3;
scale2(1462) <= r;
scale2(1463) <= d_2;
scale2(1464) <= d_2;
scale2(1465) <= d_2;
scale2(1466) <= r;
scale2(1467) <= d_3;
scale2(1468) <= d_3;
scale2(1469) <= d_3;
scale2(1470) <= r;
scale2(1471) <= d_2;
scale2(1472) <= d_2;
scale2(1473) <= d_2;
scale2(1474) <= r;
scale2(1475) <= d_3;
scale2(1476) <= d_3;
scale2(1477) <= d_3;
scale2(1478) <= r;
scale2(1479) <= d_2;
scale2(1480) <= d_2;
scale2(1481) <= d_2;
scale2(1482) <= r;
scale2(1483) <= d_3;
scale2(1484) <= d_3;
scale2(1485) <= d_3;
scale2(1486) <= r;
------------------47
scale2(1487) <= c_2;
scale2(1488) <= c_2;
scale2(1489) <= c_2;
scale2(1490) <= r;
scale2(1491) <= c_3;
scale2(1492) <= c_3;
scale2(1493) <= c_3;
scale2(1494) <= r;
scale2(1495) <= c_2;
scale2(1496) <= c_2;
scale2(1497) <= c_2;
scale2(1498) <= r;
scale2(1499) <= c_3;
scale2(1500) <= c_3;
scale2(1501) <= c_3;
scale2(1502) <= r;
scale2(1503) <= f_1;
scale2(1504) <= f_1;
scale2(1505) <= f_1;
scale2(1506) <= r;
scale2(1507) <= c_2;
scale2(1508) <= c_2;
scale2(1509) <= c_2;
scale2(1510) <= r;
scale2(1511) <= f_1;
scale2(1512) <= f_1;
scale2(1513) <= f_1;
scale2(1514) <= r;
scale2(1515) <= c_2;
scale2(1516) <= c_2;
scale2(1517) <= c_2;
scale2(1518) <= r;
------------------48
scale2(1519) <= bm_2;
scale2(1520) <= bm_2;
scale2(1521) <= bm_2;
scale2(1522) <= bm_2;
scale2(1523) <= bm_2;
scale2(1524) <= bm_2;
scale2(1525) <= bm_2;
scale2(1526) <= bm_2;
scale2(1527) <= bm_2;
scale2(1528) <= bm_2;
scale2(1529) <= bm_2;
scale2(1530) <= bm_2;
scale2(1531) <= bm_2;
scale2(1532) <= bm_2;
scale2(1533) <= bm_2;
scale2(1534) <= bm_2;
scale2(1535) <= bm_2;
scale2(1536) <= bm_2;
scale2(1537) <= bm_2;
scale2(1538) <= r;
scale2(1539) <= f_1;
scale2(1540) <= f_1;
scale2(1541) <= f_1;
scale2(1542) <= r;
scale2(1543) <= g_1;
scale2(1544) <= g_1;
scale2(1545) <= g_1;
scale2(1546) <= r;
scale2(1547) <= a_2;
scale2(1548) <= a_2;
scale2(1549) <= a_2;
scale2(1550) <= a_2;



		

process (n_clk,rss,rst)
begin
   if rss = '1' or rst = '1' then
      dot_data_00 <= zr;
		dot_data_01 <= zr;
		dot_data_02 <= zr;
		dot_data_03 <= zr;
		dot_data_04 <= zr;
		dot_data_05 <= zr;
		dot_data_06 <= zr;
		dot_data_07 <= zr;
		dot_data_08 <= zr;
		dot_data_09 <= zr;
		dot_data_10 <= zr;
		dot_data_11 <= zr;
		dot_data_12 <= zr;
		dot_data_13 <= zr;
		d_dp <= zr;
		d_d  <= zr;
		d_dm <= zr;		
	elsif n_clk'event and n_clk = '1' then
		d_dp        <= dot_data_00;
		d_d         <= dot_data_01;
		d_dm        <= dot_data_02;
		dot_data_00 <= dot_data_01;
		dot_data_01 <= dot_data_02;
		dot_data_02 <= dot_data_03;
		dot_data_03 <= dot_data_04;
		dot_data_04 <= dot_data_05;
		dot_data_05 <= dot_data_06;
		dot_data_06 <= dot_data_07;
		dot_data_07 <= dot_data_08;
		dot_data_08 <= dot_data_09;
		dot_data_09 <= dot_data_10;
		dot_data_10 <= dot_data_11;
		dot_data_11 <= dot_data_12;
		dot_data_12 <= dot_data_13;
		dot_data_13 <= data_b(note);
	end if;
end process;




u0 : dot_dis
port map (
	clk => clk,
	dot_data_00 => dot_data_00,
	dot_data_01 => dot_data_01,
	dot_data_02 => dot_data_02,
	dot_data_03 => dot_data_03,
	dot_data_04 => dot_data_04,
	dot_data_05 => dot_data_05,
	dot_data_06 => dot_data_06,
	dot_data_07 => dot_data_07,
	dot_data_08 => dot_data_08,
	dot_data_09 => dot_data_09,
	dot_data_10 => dot_data_10,
	dot_data_11 => dot_data_11,
	dot_data_12 => dot_data_12,
	dot_data_13 => dot_data_13,
	dot_d => dot_d,
	dot_scan => dot_scan 
);
----------------------------------------------------------------piezo
-------------dot + 15
scale(0) <= r;
scale(1) <= r;
scale(2) <= r;
scale(3) <= r;
scale(4) <= r;
scale(5) <= r;
scale(6) <= r;
scale(7) <= r;
scale(8) <= r;
scale(9) <= r;
scale(10) <= r;
scale(11) <= r;
scale(12) <= r;
scale(13) <= r;
scale(14) <= r;
------------------1
scale(15) <= bm_5;
scale(16) <= bm_5;
scale(17) <= bm_5;
scale(18) <= r;
scale(19) <= a_5;
scale(20) <= a_5;
scale(21) <= a_5;
scale(22) <= r;
scale(23) <= g_4;
scale(24) <= g_4;
scale(25) <= g_4;
scale(26) <= g_4;
scale(27) <= g_4;
scale(28) <= r;
scale(29) <= f_4;
scale(30) <= r;
scale(31) <= a_5;
scale(32) <= a_5;
scale(33) <= a_5;
scale(34) <= r;
scale(35) <= g_4;
scale(36) <= g_4;
scale(37) <= g_4;
scale(38) <= r;
scale(39) <= f_4;
scale(40) <= f_4;
scale(41) <= f_4;
scale(42) <= r;
scale(43) <= em_4;
scale(44) <= em_4;
scale(45) <= em_4;
scale(46) <= r;
-----------------------2
scale(47) <= g_4;
scale(48) <= g_4;
scale(49) <= g_4;
scale(50) <= r;
scale(51) <= f_4;
scale(52) <= f_4;
scale(53) <= f_4;
scale(54) <= r;
scale(55) <= em_4;
scale(56) <= r;
scale(57) <= d_4;
scale(58) <= d_4;
scale(59) <= d_4;
scale(60) <= d_4;
scale(61) <= d_4;
scale(62) <= r;
scale(63) <= f_4;
scale(64) <= f_4;
scale(65) <= f_4;
scale(66) <= f_4;
scale(67) <= f_4;
scale(68) <= f_4;
scale(69) <= f_4;
scale(70) <= f_4;
scale(71) <= f_4;
scale(72) <= f_4;
scale(73) <= f_4;
scale(74) <= r;
scale(75) <= d_4;
scale(76) <= r;
scale(77) <= c_4;
scale(78) <= r;
---------------------3
scale(79) <= bm_4;
scale(80) <= bm_4;
scale(81) <= bm_4;
scale(82) <= r;
scale(83) <= c_4;
scale(84) <= c_4;
scale(85) <= c_4;
scale(86) <= r;
scale(87) <= d_4;
scale(88) <= d_4;
scale(89) <= d_4;
scale(90) <= r;
scale(91) <= em_4;
scale(92) <= em_4;
scale(93) <= em_4;
scale(94) <= r;
scale(95) <= c_4;
scale(96) <= c_4;
scale(97) <= c_4;
scale(98) <= r;
scale(99) <= d_4;
scale(100) <= r;
scale(101) <= em_4;
scale(102) <= em_4;
scale(103) <= em_4;
scale(104) <= em_4;
scale(105) <= em_4;
scale(106) <= r;
scale(107) <= f_4;
scale(108) <= f_4;
scale(109) <= f_4;
scale(110) <= r;
-------------------4
scale(111) <= f_4;
scale(112) <= f_4;
scale(113) <= f_4;
scale(114) <= r;
scale(115) <= g_4;
scale(116) <= g_4;
scale(117) <= g_4;
scale(118) <= r;
scale(119) <= a_5;
scale(120) <= r;
scale(121) <= g_4;
scale(122) <= g_4;
scale(123) <= g_4;
scale(124) <= g_4;
scale(125) <= g_4;
scale(126) <= r;
scale(127) <= f_4;
scale(128) <= f_4;
scale(129) <= f_4;
scale(130) <= r;
scale(131) <= f_4;
scale(132) <= f_4;
scale(133) <= f_4;
scale(134) <= r;
scale(135) <= g_4;
scale(136) <= g_4;
scale(137) <= g_4;
scale(138) <= r;
scale(139) <= a_5;
scale(140) <= a_5;
scale(141) <= a_5;
scale(142) <= r;
------------------5
scale(143) <= bm_5;
scale(144) <= bm_5;
scale(145) <= bm_5;
scale(146) <= r;
scale(147) <= a_5;
scale(148) <= a_5;
scale(149) <= a_5;
scale(150) <= r;
scale(151) <= g_4;
scale(152) <= g_4;
scale(153) <= g_4;
scale(154) <= g_4;
scale(155) <= g_4;
scale(156) <= r;
scale(157) <= f_4;
scale(158) <= r;
scale(159) <= a_5;
scale(160) <= a_5;
scale(161) <= a_5;
scale(162) <= r;
scale(163) <= g_4;
scale(164) <= g_4;
scale(165) <= g_4;
scale(166) <= r;
scale(167) <= f_4;
scale(168) <= f_4;
scale(169) <= f_4;
scale(170) <= r;
scale(171) <= em_4;
scale(172) <= em_4;
scale(173) <= em_4;
scale(174) <= r;
-----------------------6
scale(175) <= g_4;
scale(176) <= g_4;
scale(177) <= g_4;
scale(178) <= r;
scale(179) <= f_4;
scale(180) <= f_4;
scale(181) <= f_4;
scale(182) <= r;
scale(183) <= em_4;
scale(184) <= r;
scale(185) <= d_4;
scale(186) <= d_4;
scale(187) <= d_4;
scale(188) <= d_4;
scale(189) <= d_4;
scale(190) <= r;
scale(191) <= f_4;
scale(192) <= f_4;
scale(193) <= f_4;
scale(194) <= f_4;
scale(195) <= f_4;
scale(196) <= f_4;
scale(197) <= f_4;
scale(198) <= f_4;
scale(199) <= f_4;
scale(200) <= f_4;
scale(201) <= f_4;
scale(202) <= r;
scale(203) <= d_4;
scale(204) <= r;
scale(205) <= c_4;
scale(206) <= r;
---------------------7
scale(207) <= bm_4;
scale(208) <= bm_4;
scale(209) <= bm_4;
scale(210) <= r;
scale(211) <= c_4;
scale(212) <= c_4;
scale(213) <= c_4;
scale(214) <= r;
scale(215) <= d_4;
scale(216) <= d_4;
scale(217) <= d_4;
scale(218) <= r;
scale(219) <= em_4;
scale(220) <= em_4;
scale(221) <= em_4;
scale(222) <= r;
scale(223) <= c_4;
scale(224) <= c_4;
scale(225) <= c_4;
scale(226) <= r;
scale(227) <= d_4;
scale(228) <= r;
scale(229) <= em_4;
scale(230) <= em_4;
scale(231) <= em_4;
scale(232) <= em_4;
scale(233) <= em_4;
scale(234) <= r;
scale(235) <= f_4;
scale(236) <= f_4;
scale(237) <= f_4;
scale(238) <= r;
---------------------------8
scale(239) <= f_4;
scale(240) <= f_4;
scale(241) <= f_4;
scale(242) <= r;
scale(243) <= g_4;
scale(244) <= g_4;
scale(245) <= g_4;
scale(246) <= r;
scale(247) <= a_5;
scale(248) <= r;
scale(249) <= f_4;
scale(250) <= f_4;
scale(251) <= f_4;
scale(252) <= f_4;
scale(253) <= f_4;
scale(254) <= r;
scale(255) <= bm_5;
scale(256) <= bm_5;
scale(257) <= bm_5;
scale(258) <= r;
scale(259) <= f_4;
scale(260) <= f_4;
scale(261) <= f_4;
scale(262) <= r;
scale(263) <= g_4;
scale(264) <= g_4;
scale(265) <= g_4;
scale(266) <= r;
scale(267) <= am_4;
scale(268) <= am_4;
scale(269) <= am_4;
scale(270) <= r;
---------------------------9
scale(271) <= a_5;
scale(272) <= a_5;
scale(273) <= a_5;
scale(274) <= a_5;
scale(275) <= f_5;
scale(276) <= f_5;
scale(277) <= f_5;
scale(278) <= r;
scale(279) <= g_5;
scale(280) <= g_5;
scale(281) <= g_5;
scale(282) <= r;
scale(283) <= am_5;
scale(284) <= am_5;
scale(285) <= am_5;
scale(286) <= r;
scale(287) <= a_6;
scale(288) <= a_6;
scale(289) <= a_6;
scale(290) <= a_6;
scale(291) <= f_4;
scale(292) <= f_4;
scale(293) <= f_4;
scale(294) <= r;
scale(295) <= g_4;
scale(296) <= g_4;
scale(297) <= g_4;
scale(298) <= r;
scale(299) <= a_5;
scale(300) <= a_5;
scale(301) <= a_5;
scale(302) <= r;
----------------------10
scale(303) <= bm_5;
scale(304) <= bm_5;
scale(305) <= bm_5;
scale(306) <= bm_5;
scale(307) <= f_5;
scale(308) <= f_5;
scale(309) <= f_5;
scale(310) <= r;
scale(311) <= g_5;
scale(312) <= g_5;
scale(313) <= g_5;
scale(314) <= r;
scale(315) <= a_6;
scale(316) <= a_6;
scale(317) <= a_6;
scale(318) <= r;
scale(319) <= bm_6;
scale(320) <= bm_6;
scale(321) <= bm_6;
scale(322) <= bm_6;
scale(323) <= f_4;
scale(324) <= f_4;
scale(325) <= f_4;
scale(326) <= r;
scale(327) <= g_4;
scale(328) <= g_4;
scale(329) <= g_4;
scale(330) <= r;
scale(331) <= a_5;
scale(332) <= a_5;
scale(333) <= a_5;
scale(334) <= r;
-----------------------------11
scale(335) <= c_5;
scale(336) <= c_5;
scale(337) <= c_5;
scale(338) <= c_5;
scale(339) <= f_5;
scale(340) <= f_5;
scale(341) <= f_5;
scale(342) <= r;
scale(343) <= g_5;
scale(344) <= g_5;
scale(345) <= g_5;
scale(346) <= r;
scale(347) <= a_6;
scale(348) <= a_6;
scale(349) <= a_6;
scale(350) <= r;
scale(351) <= c_6;
scale(352) <= c_6;
scale(353) <= c_6;
scale(354) <= c_6;
scale(355) <= f_4;
scale(356) <= f_4;
scale(357) <= f_4;
scale(358) <= r; 
scale(359) <= g_4;
scale(360) <= g_4;
scale(361) <= g_4;
scale(362) <= r;
scale(363) <= a_5;
scale(364) <= a_5;
scale(365) <= a_5;
scale(366) <= r;
----------------------------12
scale(367) <= d_5;
scale(368) <= d_5;
scale(369) <= d_5;
scale(370) <= d_5;
scale(371) <= f_5;
scale(372) <= f_5;
scale(373) <= f_5;
scale(374) <= r;
scale(375) <= g_5;
scale(376) <= g_5;
scale(377) <= g_5;
scale(378) <= r;
scale(379) <= a_6;
scale(380) <= a_6;
scale(381) <= a_6;
scale(382) <= r;
scale(383) <= d_6;
scale(384) <= d_6;
scale(385) <= d_6;
scale(386) <= d_6;
scale(387) <= bm_5;
scale(388) <= bm_5;
scale(389) <= bm_5;
scale(390) <= r;
scale(391) <= c_5;
scale(392) <= c_5;
scale(393) <= c_5;
scale(394) <= r;
scale(395) <= d_5;
scale(396) <= d_5; 
scale(397) <= d_5;
scale(398) <= r;
--------------------13
scale(399) <= em_5;
scale(400) <= em_5;
scale(401) <= em_5;
scale(402) <= r;
scale(403) <= em_5;
scale(404) <= em_5;
scale(405) <= em_5;
scale(406) <= em_5;
scale(407) <= em_5;
scale(408) <= em_5;
scale(409) <= em_5;
scale(410) <= r; 
scale(411) <= em_5;
scale(412) <= em_5;
scale(413) <= em_5;
scale(414) <= em_5;
scale(415) <= em_5;
scale(416) <= em_5;
scale(417) <= em_5;
scale(418) <= r;
scale(419) <= d_5;
scale(420) <= d_5;
scale(421) <= d_5;
scale(422) <= r;
scale(423) <= c_5;
scale(424) <= c_5;
scale(425) <= c_5;
scale(426) <= c_5;
scale(427) <= c_5;
scale(428) <= c_5;
scale(429) <= c_5;
scale(430) <= r;
----------------------14
scale(431) <= d_5;
scale(432) <= d_5;
scale(433) <= d_5;
scale(434) <= d_5;
scale(435) <= d_5;
scale(436) <= d_5;
scale(437) <= d_5;
scale(438) <= d_5;
scale(439) <= d_5;
scale(440) <= d_5;
scale(441) <= d_5;
scale(442) <= d_5;
scale(443) <= d_5;
scale(444) <= d_5; 
scale(445) <= d_5;
scale(446) <= d_5;
scale(447) <= d_5;
scale(448) <= d_5;
scale(449) <= d_5;
scale(450) <= d_5;
scale(451) <= d_5;
scale(452) <= d_5;
scale(453) <= d_5;
scale(454) <= r;
scale(455) <= d_5;
scale(456) <= d_5;
scale(457) <= d_5;
scale(458) <= d_5;
scale(459) <= d_5;
scale(460) <= d_5;
scale(461) <= d_5;
scale(462) <= r;
-----------------------15
scale(463) <= c_5;
scale(464) <= c_5;
scale(465) <= c_5;
scale(466) <= c_5;
scale(467) <= c_5;
scale(468) <= c_5;
scale(469) <= c_5;
scale(470) <= c_5;
scale(471) <= c_5;
scale(472) <= c_5;
scale(473) <= c_5;
scale(474) <= r;
scale(475) <= g_4;
scale(476) <= g_4;
scale(477) <= g_4;
scale(478) <= g_4;
scale(479) <= g_4;
scale(480) <= g_4;
scale(481) <= g_4;
scale(482) <= r;
scale(483) <= g_4;
scale(484) <= g_4;
scale(485) <= g_4;
scale(486) <= r;
scale(487) <= d_5;
scale(488) <= d_5;
scale(489) <= d_5;
scale(490) <= d_5;
scale(491) <= d_5;
scale(492) <= d_5;
scale(493) <= d_5;
scale(494) <= r;
------------------16
scale(495) <= c_5;
scale(496) <= c_5;
scale(497) <= c_5;
scale(498) <= c_5;
scale(499) <= c_5;
scale(500) <= c_5;
scale(501) <= c_5;
scale(502) <= c_5;
scale(503) <= c_5;
scale(504) <= c_5;
scale(505) <= c_5;
scale(506) <= c_5;
scale(507) <= c_5;
scale(508) <= c_5;
scale(509) <= c_5;
scale(510) <= c_5;
scale(511) <= c_5;
scale(512) <= c_5;
scale(513) <= c_5;
scale(514) <= r;
scale(515) <= f_4;
scale(516) <= f_4;
scale(517) <= f_4;
scale(518) <= r;
scale(519) <= g_4;
scale(520) <= g_4;
scale(521) <= g_4;
scale(522) <= r;
scale(523) <= am_4;
scale(524) <= am_4;
scale(525) <= am_4;
scale(526) <= r;
---------------------------17
scale(527) <= a_5;
scale(528) <= a_5;
scale(529) <= a_5;
scale(530) <= a_5;
scale(531) <= f_5;
scale(532) <= f_5;
scale(533) <= f_5;
scale(534) <= r;
scale(535) <= g_5;
scale(536) <= g_5;
scale(537) <= g_5;
scale(538) <= r;
scale(539) <= am_5;
scale(540) <= am_5;
scale(541) <= am_5;
scale(542) <= r;
scale(543) <= a_6;
scale(544) <= a_6;
scale(545) <= a_6;
scale(546) <= a_6;
scale(547) <= f_4;
scale(548) <= f_4;
scale(549) <= f_4;
scale(550) <= r;
scale(551) <= g_4;
scale(552) <= g_4;
scale(553) <= g_4;
scale(554) <= r;
scale(555) <= a_5;
scale(556) <= a_5;
scale(557) <= a_5;
scale(558) <= r;
----------------------18
scale(559) <= bm_5;
scale(560) <= bm_5;
scale(561) <= bm_5;
scale(562) <= bm_5;
scale(563) <= f_5;
scale(564) <= f_5;
scale(565) <= f_5;
scale(566) <= r;
scale(567) <= g_5;
scale(568) <= g_5;
scale(569) <= g_5;
scale(570) <= r;
scale(571) <= a_6;
scale(572) <= a_6;
scale(573) <= a_6;
scale(574) <= r;
scale(575) <= bm_6;
scale(576) <= bm_6;
scale(577) <= bm_6;
scale(578) <= bm_6;
scale(579) <= f_4;
scale(580) <= f_4;
scale(581) <= f_4;
scale(582) <= r;
scale(583) <= g_4;
scale(584) <= g_4;
scale(585) <= g_4;
scale(586) <= r;
scale(587) <= a_5;
scale(588) <= a_5;
scale(589) <= a_5;
scale(590) <= r;
-----------------------------19
scale(591) <= c_5;
scale(592) <= c_5;
scale(593) <= c_5;
scale(594) <= c_5;
scale(595) <= f_5;
scale(596) <= f_5;
scale(597) <= f_5;
scale(598) <= r;
scale(599) <= g_5;
scale(600) <= g_5;
scale(601) <= g_5;
scale(602) <= r;
scale(603) <= a_6;
scale(604) <= a_6;
scale(605) <= a_6;
scale(606) <= r;
scale(607) <= c_6;
scale(608) <= c_6;
scale(609) <= c_6;
scale(610) <= c_6;
scale(611) <= f_4;
scale(612) <= f_4;
scale(613) <= f_4;
scale(614) <= r; 
scale(615) <= g_4;
scale(616) <= g_4;
scale(617) <= g_4;
scale(618) <= r;
scale(619) <= a_5;
scale(620) <= a_5;
scale(621) <= a_5;
scale(622) <= r;
----------------------------20
scale(623) <= d_5;
scale(624) <= d_5;
scale(625) <= d_5;
scale(626) <= d_5;
scale(627) <= f_5;
scale(628) <= f_5;
scale(629) <= f_5;
scale(630) <= r;
scale(631) <= g_5;
scale(632) <= g_5;
scale(633) <= g_5;
scale(634) <= r;
scale(635) <= a_6;
scale(636) <= a_6;
scale(637) <= a_6;
scale(638) <= r;
scale(639) <= d_6;
scale(640) <= d_6;
scale(641) <= d_6;
scale(642) <= d_6;
scale(643) <= bm_5;
scale(644) <= bm_5;
scale(645) <= bm_5;
scale(646) <= r;
scale(647) <= c_5;
scale(648) <= c_5;
scale(649) <= c_5;
scale(650) <= r;
scale(651) <= d_5;
scale(652) <= d_5; 
scale(653) <= d_5;
scale(654) <= r;
--------------------------------21
scale(655) <= em_5;
scale(656) <= em_5;
scale(657) <= em_5;
scale(658) <= r;
scale(659) <= em_5;
scale(660) <= em_5;
scale(661) <= em_5;
scale(662) <= em_5;
scale(663) <= em_5;
scale(664) <= em_5;
scale(665) <= em_5;
scale(666) <= r; 
scale(667) <= em_5;
scale(668) <= em_5;
scale(669) <= em_5;
scale(670) <= em_5;
scale(671) <= em_5;
scale(672) <= em_5;
scale(673) <= em_5;
scale(674) <= r;
scale(675) <= d_5;
scale(676) <= d_5;
scale(677) <= d_5;
scale(678) <= r;
scale(679) <= c_5;
scale(680) <= c_5;
scale(681) <= c_5;
scale(682) <= c_5;
scale(683) <= c_5;
scale(684) <= c_5;
scale(685) <= c_5;
scale(686) <= r;
----------------------22
scale(687) <= d_5;
scale(688) <= d_5;
scale(689) <= d_5;
scale(690) <= d_5;
scale(691) <= d_5;
scale(692) <= d_5;
scale(693) <= d_5;
scale(694) <= d_5;
scale(695) <= d_5;
scale(696) <= d_5;
scale(697) <= d_5;
scale(698) <= d_5;
scale(699) <= d_5;
scale(700) <= d_5; 
scale(701) <= d_5;
scale(702) <= d_5;
scale(703) <= d_5;
scale(704) <= d_5;
scale(705) <= d_5;
scale(706) <= d_5;
scale(707) <= d_5;
scale(708) <= d_5;
scale(709) <= d_5;
scale(710) <= r;
scale(711) <= d_5;
scale(712) <= d_5;
scale(713) <= d_5;
scale(714) <= d_5;
scale(715) <= d_5;
scale(716) <= d_5;
scale(717) <= d_5;
scale(718) <= r;
-------------------23
scale(719) <= c_5;
scale(720) <= c_5;
scale(721) <= c_5;
scale(722) <= c_5;
scale(723) <= c_5;
scale(724) <= c_5;
scale(725) <= c_5;
scale(726) <= c_5;
scale(727) <= c_5;
scale(728) <= c_5;
scale(729) <= c_5;
scale(730) <= r;
scale(731) <= f_4;
scale(732) <= f_4;
scale(733) <= f_4;
scale(734) <= f_4;
scale(735) <= f_4;
scale(736) <= f_4;
scale(737) <= f_4;
scale(738) <= r; 
scale(739) <= d_5;
scale(740) <= d_5;
scale(741) <= d_5;
scale(742) <= r;
scale(743) <= f_4;
scale(744) <= f_4;
scale(745) <= f_4;
scale(746) <= r;
scale(747) <= d_5;
scale(748) <= d_5;
scale(749) <= d_5;
scale(750) <= r;
----------------------------------24
scale(751) <= bm_5;
scale(752) <= bm_5;
scale(753) <= bm_5;
scale(754) <= bm_5;
scale(755) <= bm_5;
scale(756) <= bm_5;
scale(757) <= bm_5;
scale(758) <= bm_5;
scale(759) <= bm_5;
scale(760) <= bm_5;
scale(761) <= bm_5;
scale(762) <= bm_5;
scale(763) <= bm_5;
scale(764) <= bm_5;
scale(765) <= bm_5;
scale(766) <= bm_5;
scale(767) <= bm_5;
scale(768) <= bm_5;
scale(769) <= bm_5;
scale(770) <= r;
scale(771) <= f_4;
scale(772) <= f_4;
scale(773) <= f_4;
scale(774) <= r;
scale(775) <= g_4;
scale(776) <= g_4;
scale(777) <= g_4;
scale(778) <= r;
scale(779) <= a_5;
scale(780) <= a_5;
scale(781) <= a_5;
scale(782) <= r;
------------------25
scale(783) <= bm_5;
scale(784) <= bm_5;
scale(785) <= bm_5;
scale(786) <= r;
scale(787) <= a_5;
scale(788) <= a_5;
scale(789) <= a_5;
scale(790) <= r;
scale(791) <= g_4;
scale(792) <= g_4;
scale(793) <= g_4;
scale(794) <= g_4;
scale(795) <= g_4;
scale(796) <= r;
scale(797) <= f_4;
scale(798) <= r;
scale(799) <= a_5;
scale(800) <= a_5;
scale(801) <= a_5;
scale(802) <= r;
scale(803) <= g_4;
scale(804) <= g_4;
scale(805) <= g_4;
scale(806) <= r;
scale(807) <= f_4;
scale(808) <= f_4;
scale(809) <= f_4;
scale(810) <= r;
scale(811) <= em_4;
scale(812) <= em_4;
scale(813) <= em_4;
scale(814) <= r;
-----------------------26
scale(815) <= g_4;
scale(816) <= g_4;
scale(817) <= g_4;
scale(818) <= r;
scale(819) <= f_4;
scale(820) <= f_4;
scale(821) <= f_4;
scale(822) <= r;
scale(823) <= em_4;
scale(824) <= r;
scale(825) <= d_4;
scale(826) <= d_4;
scale(827) <= d_4;
scale(828) <= d_4;
scale(829) <= d_4;
scale(830) <= r;
scale(831) <= f_4;
scale(832) <= f_4;
scale(833) <= f_4;
scale(834) <= f_4;
scale(835) <= f_4;
scale(836) <= f_4;
scale(837) <= f_4;
scale(838) <= f_4;
scale(839) <= f_4;
scale(840) <= f_4;
scale(841) <= f_4;
scale(842) <= r;
scale(843) <= d_4;
scale(844) <= r;
scale(845) <= c_4;
scale(846) <= r;
---------------------27
scale(847) <= bm_4;
scale(848) <= bm_4;
scale(849) <= bm_4;
scale(850) <= r;
scale(851) <= c_4;
scale(852) <= c_4;
scale(853) <= c_4;
scale(854) <= r;
scale(855) <= d_4;
scale(856) <= d_4;
scale(857) <= d_4;
scale(858) <= r;
scale(859) <= em_4;
scale(860) <= em_4;
scale(861) <= em_4;
scale(862) <= r;
scale(863) <= c_4;
scale(864) <= c_4;
scale(865) <= c_4;
scale(866) <= r;
scale(867) <= d_4;
scale(868) <= r;
scale(869) <= em_4;
scale(870) <= em_4;
scale(871) <= em_4;
scale(872) <= em_4;
scale(873) <= em_4;
scale(874) <= r;
scale(875) <= f_4;
scale(876) <= f_4;
scale(877) <= f_4;
scale(878) <= r;
-------------------28
scale(879) <= f_4;
scale(880) <= f_4;
scale(881) <= f_4;
scale(882) <= r;
scale(883) <= g_4;
scale(884) <= g_4;
scale(885) <= g_4;
scale(886) <= r;
scale(887) <= a_5;
scale(888) <= r;
scale(889) <= g_4;
scale(890) <= g_4;
scale(891) <= g_4;
scale(892) <= g_4;
scale(893) <= g_4;
scale(894) <= r;
scale(895) <= f_4;
scale(896) <= f_4;
scale(897) <= f_4;
scale(898) <= r;
scale(899) <= f_4;
scale(900) <= f_4;
scale(901) <= f_4;
scale(902) <= r;
scale(903) <= g_4;
scale(904) <= g_4;
scale(905) <= g_4;
scale(906) <= r;
scale(907) <= a_5;
scale(908) <= a_5;
scale(909) <= a_5;
scale(910) <= r;
------------------29
scale(911) <= bm_5;
scale(912) <= bm_5;
scale(913) <= bm_5;
scale(914) <= r;
scale(915) <= a_5;
scale(916) <= a_5;
scale(917) <= a_5;
scale(918) <= r;
scale(919) <= g_4;
scale(920) <= g_4;
scale(921) <= g_4;
scale(922) <= g_4;
scale(923) <= g_4;
scale(924) <= r;
scale(925) <= f_4;
scale(926) <= r;
scale(927) <= a_5;
scale(928) <= a_5;
scale(929) <= a_5;
scale(930) <= r;
scale(931) <= g_4;
scale(932) <= g_4;
scale(933) <= g_4;
scale(934) <= r;
scale(935) <= f_4;
scale(936) <= f_4;
scale(937) <= f_4;
scale(938) <= r;
scale(939) <= em_4;
scale(940) <= em_4;
scale(941) <= em_4;
scale(942) <= r;
-----------------------30
scale(943) <= g_4;
scale(944) <= g_4;
scale(945) <= g_4;
scale(946) <= r;
scale(947) <= f_4;
scale(948) <= f_4;
scale(949) <= f_4;
scale(950) <= r;
scale(951) <= em_4;
scale(952) <= r;
scale(953) <= d_4;
scale(954) <= d_4;
scale(955) <= d_4;
scale(956) <= d_4;
scale(957) <= d_4;
scale(958) <= r;
scale(959) <= f_4;
scale(960) <= f_4;
scale(961) <= f_4;
scale(962) <= f_4;
scale(963) <= f_4;
scale(964) <= f_4;
scale(965) <= f_4;
scale(966) <= f_4;
scale(967) <= f_4;
scale(968) <= f_4;
scale(969) <= f_4;
scale(970) <= r;
scale(971) <= d_4;
scale(972) <= r;
scale(973) <= c_4;
scale(974) <= r;
---------------------31
scale(975) <= bm_4;
scale(976) <= bm_4;
scale(977) <= bm_4;
scale(978) <= r;
scale(979) <= c_4;
scale(980) <= c_4;
scale(981) <= c_4;
scale(982) <= r;
scale(983) <= d_4;
scale(984) <= d_4;
scale(985) <= d_4;
scale(986) <= r;
scale(987) <= em_4;
scale(988) <= em_4;
scale(989) <= em_4;
scale(990) <= r;
scale(991) <= c_4;
scale(992) <= c_4;
scale(993) <= c_4;
scale(994) <= r;
scale(995) <= d_4;
scale(996) <= r;
scale(997) <= em_4;
scale(998) <= em_4;
scale(999) <= em_4;
scale(1000) <= em_4;
scale(1001) <= em_4;
scale(1002) <= r;
scale(1003) <= f_4;
scale(1004) <= f_4;
scale(1005) <= f_4;
scale(1006) <= r;
---------------------------32
scale(1007) <= f_4;
scale(1008) <= f_4;
scale(1009) <= f_4;
scale(1010) <= r;
scale(1011) <= g_4;
scale(1012) <= g_4;
scale(1013) <= g_4;
scale(1014) <= r;
scale(1015) <= a_5;
scale(1016) <= r;
scale(1017) <= f_4;
scale(1018) <= f_4;
scale(1019) <= f_4;
scale(1020) <= f_4;
scale(1021) <= f_4;
scale(1022) <= r;
scale(1023) <= bm_5;
scale(1024) <= bm_5;
scale(1025) <= bm_5;
scale(1026) <= r;
scale(1027) <= f_4;
scale(1028) <= f_4;
scale(1029) <= f_4;
scale(1030) <= r;
scale(1031) <= g_4;
scale(1032) <= g_4;
scale(1033) <= g_4;
scale(1034) <= r;
scale(1035) <= am_4;
scale(1036) <= am_4;
scale(1037) <= am_4;
scale(1038) <= r;
---------------------------33
scale(1039) <= a_5;
scale(1040) <= a_5;
scale(1041) <= a_5;
scale(1042) <= a_5;
scale(1043) <= f_5;
scale(1044) <= f_5;
scale(1045) <= f_5;
scale(1046) <= r;
scale(1047) <= g_5;
scale(1048) <= g_5;
scale(1049) <= g_5;
scale(1050) <= r;
scale(1051) <= am_5;
scale(1052) <= am_5;
scale(1053) <= am_5;
scale(1054) <= r;
scale(1055) <= a_6;
scale(1056) <= a_6;
scale(1057) <= a_6;
scale(1058) <= a_6;
scale(1059) <= f_4;
scale(1060) <= f_4;
scale(1061) <= f_4;
scale(1062) <= r;
scale(1063) <= g_4;
scale(1064) <= g_4;
scale(1065) <= g_4;
scale(1066) <= r;
scale(1067) <= a_5;
scale(1068) <= a_5;
scale(1069) <= a_5;
scale(1070) <= r;
----------------------34
scale(1071) <= bm_5;
scale(1072) <= bm_5;
scale(1073) <= bm_5;
scale(1074) <= bm_5;
scale(1075) <= f_5;
scale(1076) <= f_5;
scale(1077) <= f_5;
scale(1078) <= r;
scale(1079) <= g_5;
scale(1080) <= g_5;
scale(1081) <= g_5;
scale(1082) <= r;
scale(1083) <= a_6;
scale(1084) <= a_6;
scale(1085) <= a_6;
scale(1086) <= r;
scale(1087) <= bm_6;
scale(1088) <= bm_6;
scale(1089) <= bm_6;
scale(1090) <= bm_6;
scale(1091) <= f_4;
scale(1092) <= f_4;
scale(1093) <= f_4;
scale(1094) <= r;
scale(1095) <= g_4;
scale(1096) <= g_4;
scale(1097) <= g_4;
scale(1098) <= r;
scale(1099) <= a_5;
scale(1100) <= a_5;
scale(1101) <= a_5;
scale(1102) <= r;
-----------------------------35
scale(1103) <= c_5;
scale(1104) <= c_5;
scale(1105) <= c_5;
scale(1106) <= c_5;
scale(1107) <= f_5;
scale(1108) <= f_5;
scale(1109) <= f_5;
scale(1110) <= r;
scale(1111) <= g_5;
scale(1112) <= g_5;
scale(1113) <= g_5;
scale(1114) <= r;
scale(1115) <= a_6;
scale(1116) <= a_6;
scale(1117) <= a_6;
scale(1118) <= r;
scale(1119) <= c_6;
scale(1120) <= c_6;
scale(1121) <= c_6;
scale(1122) <= c_6;
scale(1123) <= f_4;
scale(1124) <= f_4;
scale(1125) <= f_4;
scale(1126) <= r; 
scale(1127) <= g_4;
scale(1128) <= g_4;
scale(1129) <= g_4;
scale(1130) <= r;
scale(1131) <= a_5;
scale(1132) <= a_5;
scale(1133) <= a_5;
scale(1134) <= r;
----------------------------36
scale(1135) <= d_5;
scale(1136) <= d_5;
scale(1137) <= d_5;
scale(1138) <= d_5;
scale(1139) <= f_5;
scale(1140) <= f_5;
scale(1141) <= f_5;
scale(1142) <= r;
scale(1143) <= g_5;
scale(1144) <= g_5;
scale(1145) <= g_5;
scale(1146) <= r;
scale(1147) <= a_6;
scale(1148) <= a_6;
scale(1149) <= a_6;
scale(1150) <= r;
scale(1151) <= d_6;
scale(1152) <= d_6;
scale(1153) <= d_6;
scale(1154) <= d_6;
scale(1155) <= bm_5;
scale(1156) <= bm_5;
scale(1157) <= bm_5;
scale(1158) <= r;
scale(1159) <= c_5;
scale(1160) <= c_5;
scale(1161) <= c_5;
scale(1162) <= r;
scale(1163) <= d_5;
scale(1164) <= d_5; 
scale(1165) <= d_5;
scale(1166) <= r;
--------------------37
scale(1167) <= em_5;
scale(1168) <= em_5;
scale(1169) <= em_5;
scale(1170) <= r;
scale(1171) <= em_5;
scale(1172) <= em_5;
scale(1173) <= em_5;
scale(1174) <= em_5;
scale(1175) <= em_5;
scale(1176) <= em_5;
scale(1177) <= em_5;
scale(1178) <= r; 
scale(1179) <= em_5;
scale(1180) <= em_5;
scale(1181) <= em_5;
scale(1182) <= em_5;
scale(1183) <= em_5;
scale(1184) <= em_5;
scale(1185) <= em_5;
scale(1186) <= r;
scale(1187) <= d_5;
scale(1188) <= d_5;
scale(1189) <= d_5;
scale(1190) <= r;
scale(1191) <= c_5;
scale(1192) <= c_5;
scale(1193) <= c_5;
scale(1194) <= c_5;
scale(1195) <= c_5;
scale(1196) <= c_5;
scale(1197) <= c_5;
scale(1198) <= r;
----------------------38
scale(1199) <= d_5;
scale(1200) <= d_5;
scale(1201) <= d_5;
scale(1202) <= d_5;
scale(1203) <= d_5;
scale(1204) <= d_5;
scale(1205) <= d_5;
scale(1206) <= d_5;
scale(1207) <= d_5;
scale(1208) <= d_5;
scale(1209) <= d_5;
scale(1210) <= d_5;
scale(1211) <= d_5;
scale(1212) <= d_5; 
scale(1213) <= d_5;
scale(1214) <= d_5;
scale(1215) <= d_5;
scale(1216) <= d_5;
scale(1217) <= d_5;
scale(1218) <= d_5;
scale(1219) <= d_5;
scale(1220) <= d_5;
scale(1221) <= d_5;
scale(1222) <= r;
scale(1223) <= d_5;
scale(1224) <= d_5;
scale(1225) <= d_5;
scale(1226) <= d_5;
scale(1227) <= d_5;
scale(1228) <= d_5;
scale(1229) <= d_5;
scale(1230) <= r;
-----------------------39
scale(1231) <= c_5;
scale(1232) <= c_5;
scale(1233) <= c_5;
scale(1234) <= c_5;
scale(1235) <= c_5;
scale(1236) <= c_5;
scale(1237) <= c_5;
scale(1238) <= c_5;
scale(1239) <= c_5;
scale(1240) <= c_5;
scale(1241) <= c_5;
scale(1242) <= r;
scale(1243) <= g_4;
scale(1244) <= g_4;
scale(1245) <= g_4;
scale(1246) <= g_4;
scale(1247) <= g_4;
scale(1248) <= g_4;
scale(1249) <= g_4;
scale(1250) <= r;
scale(1251) <= g_4;
scale(1252) <= g_4;
scale(1253) <= g_4;
scale(1254) <= r;
scale(1255) <= d_5;
scale(1256) <= d_5;
scale(1257) <= d_5;
scale(1258) <= d_5;
scale(1259) <= d_5;
scale(1260) <= d_5;
scale(1261) <= d_5;
scale(1262) <= r;
------------------40
scale(1263) <= c_5;
scale(1264) <= c_5;
scale(1265) <= c_5;
scale(1266) <= c_5;
scale(1267) <= c_5;
scale(1268) <= c_5;
scale(1269) <= c_5;
scale(1270) <= c_5;
scale(1271) <= c_5;
scale(1272) <= c_5;
scale(1273) <= c_5;
scale(1274) <= c_5;
scale(1275) <= c_5;
scale(1276) <= c_5;
scale(1277) <= c_5;
scale(1278) <= c_5;
scale(1279) <= c_5;
scale(1280) <= c_5;
scale(1281) <= c_5;
scale(1282) <= r;
scale(1283) <= f_4;
scale(1284) <= f_4;
scale(1285) <= f_4;
scale(1286) <= r;
scale(1287) <= g_4;
scale(1288) <= g_4;
scale(1289) <= g_4;
scale(1290) <= r;
scale(1291) <= am_4;
scale(1292) <= am_4;
scale(1293) <= am_4;
scale(1294) <= r;
---------------------------41
scale(1295) <= a_5;
scale(1296) <= a_5;
scale(1297) <= a_5;
scale(1298) <= a_5;
scale(1299) <= f_5;
scale(1300) <= f_5;
scale(1301) <= f_5;
scale(1302) <= r;
scale(1303) <= g_5;
scale(1304) <= g_5;
scale(1305) <= g_5;
scale(1306) <= r;
scale(1307) <= am_5;
scale(1308) <= am_5;
scale(1309) <= am_5;
scale(1310) <= r;
scale(1311) <= a_6;
scale(1312) <= a_6;
scale(1313) <= a_6;
scale(1314) <= a_6;
scale(1315) <= f_4;
scale(1316) <= f_4;
scale(1317) <= f_4;
scale(1318) <= r;
scale(1319) <= g_4;
scale(1320) <= g_4;
scale(1321) <= g_4;
scale(1322) <= r;
scale(1323) <= a_5;
scale(1324) <= a_5;
scale(1325) <= a_5;
scale(1326) <= r;
----------------------42
scale(1327) <= bm_5;
scale(1328) <= bm_5;
scale(1329) <= bm_5;
scale(1330) <= bm_5;
scale(1331) <= f_5;
scale(1332) <= f_5;
scale(1333) <= f_5;
scale(1334) <= r;
scale(1335) <= g_5;
scale(1336) <= g_5;
scale(1337) <= g_5;
scale(1338) <= r;
scale(1339) <= a_6;
scale(1340) <= a_6;
scale(1341) <= a_6;
scale(1342) <= r;
scale(1343) <= bm_6;
scale(1344) <= bm_6;
scale(1345) <= bm_6;
scale(1346) <= bm_6;
scale(1347) <= f_4;
scale(1348) <= f_4;
scale(1349) <= f_4;
scale(1350) <= r;
scale(1351) <= g_4;
scale(1352) <= g_4;
scale(1353) <= g_4;
scale(1354) <= r;
scale(1355) <= a_5;
scale(1356) <= a_5;
scale(1357) <= a_5;
scale(1358) <= r;
-----------------------------43
scale(1359) <= c_5;
scale(1360) <= c_5;
scale(1361) <= c_5;
scale(1362) <= c_5;
scale(1363) <= f_5;
scale(1364) <= f_5;
scale(1365) <= f_5;
scale(1366) <= r;
scale(1367) <= g_5;
scale(1368) <= g_5;
scale(1369) <= g_5;
scale(1370) <= r;
scale(1371) <= a_6;
scale(1372) <= a_6;
scale(1373) <= a_6;
scale(1374) <= r;
scale(1375) <= c_6;
scale(1376) <= c_6;
scale(1377) <= c_6;
scale(1378) <= c_6;
scale(1379) <= f_4;
scale(1380) <= f_4;
scale(1381) <= f_4;
scale(1382) <= r; 
scale(1383) <= g_4;
scale(1384) <= g_4;
scale(1385) <= g_4;
scale(1386) <= r;
scale(1387) <= a_5;
scale(1388) <= a_5;
scale(1389) <= a_5;
scale(1390) <= r;
----------------------------44
scale(1391) <= d_5;
scale(1392) <= d_5;
scale(1393) <= d_5;
scale(1394) <= d_5;
scale(1395) <= f_5;
scale(1396) <= f_5;
scale(1397) <= f_5;
scale(1398) <= r;
scale(1399) <= g_5;
scale(1400) <= g_5;
scale(1401) <= g_5;
scale(1402) <= r;
scale(1403) <= a_6;
scale(1404) <= a_6;
scale(1405) <= a_6;
scale(1406) <= r;
scale(1407) <= d_6;
scale(1408) <= d_6;
scale(1409) <= d_6;
scale(1410) <= d_6;
scale(1411) <= bm_5;
scale(1412) <= bm_5;
scale(1413) <= bm_5;
scale(1414) <= r;
scale(1415) <= c_5;
scale(1416) <= c_5;
scale(1417) <= c_5;
scale(1418) <= r;
scale(1419) <= d_5;
scale(1420) <= d_5; 
scale(1421) <= d_5;
scale(1422) <= r;
--------------------------------45
scale(1423) <= em_5;
scale(1424) <= em_5;
scale(1425) <= em_5;
scale(1426) <= r;
scale(1427) <= em_5;
scale(1428) <= em_5;
scale(1429) <= em_5;
scale(1430) <= em_5;
scale(1431) <= em_5;
scale(1432) <= em_5;
scale(1433) <= em_5;
scale(1434) <= r; 
scale(1435) <= em_5;
scale(1436) <= em_5;
scale(1437) <= em_5;
scale(1438) <= em_5;
scale(1439) <= em_5;
scale(1440) <= em_5;
scale(1441) <= em_5;
scale(1442) <= r;
scale(1443) <= d_5;
scale(1444) <= d_5;
scale(1445) <= d_5;
scale(1446) <= r;
scale(1447) <= c_5;
scale(1448) <= c_5;
scale(1449) <= c_5;
scale(1450) <= c_5;
scale(1451) <= c_5;
scale(1452) <= c_5;
scale(1453) <= c_5;
scale(1454) <= r;
----------------------46
scale(1455) <= d_5;
scale(1456) <= d_5;
scale(1457) <= d_5;
scale(1458) <= d_5;
scale(1459) <= d_5;
scale(1460) <= d_5;
scale(1461) <= d_5;
scale(1462) <= d_5;
scale(1463) <= d_5;
scale(1464) <= d_5;
scale(1465) <= d_5;
scale(1466) <= d_5;
scale(1467) <= d_5;
scale(1468) <= d_5; 
scale(1469) <= d_5;
scale(1470) <= d_5;
scale(1471) <= d_5;
scale(1472) <= d_5;
scale(1473) <= d_5;
scale(1474) <= d_5;
scale(1475) <= d_5;
scale(1476) <= d_5;
scale(1477) <= d_5;
scale(1478) <= r;
scale(1479) <= d_5;
scale(1480) <= d_5;
scale(1481) <= d_5;
scale(1482) <= d_5;
scale(1483) <= d_5;
scale(1484) <= d_5;
scale(1485) <= d_5;
scale(1486) <= r;
-------------------47
scale(1487) <= c_5;
scale(1488) <= c_5;
scale(1489) <= c_5;
scale(1490) <= c_5;
scale(1491) <= c_5;
scale(1492) <= c_5;
scale(1493) <= c_5;
scale(1494) <= c_5;
scale(1495) <= c_5;
scale(1496) <= c_5;
scale(1497) <= c_5;
scale(1498) <= r;
scale(1499) <= f_4;
scale(1500) <= f_4;
scale(1501) <= f_4;
scale(1502) <= f_4;
scale(1503) <= f_4;
scale(1504) <= f_4;
scale(1505) <= f_4;
scale(1506) <= r; 
scale(1507) <= d_5;
scale(1508) <= d_5;
scale(1509) <= d_5;
scale(1510) <= r;
scale(1511) <= f_4;
scale(1512) <= f_4;
scale(1513) <= f_4;
scale(1514) <= r;
scale(1515) <= d_5;
scale(1516) <= d_5;
scale(1517) <= d_5;
scale(1518) <= r;
----------------------------------48
scale(1519) <= bm_5;
scale(1520) <= bm_5;
scale(1521) <= bm_5;
scale(1522) <= bm_5;
scale(1523) <= bm_5;
scale(1524) <= bm_5;
scale(1525) <= bm_5;
scale(1526) <= bm_5;
scale(1527) <= bm_5;
scale(1528) <= bm_5;
scale(1529) <= bm_5;
scale(1530) <= bm_5;
scale(1531) <= bm_5;
scale(1532) <= bm_5;
scale(1533) <= bm_5;
scale(1534) <= bm_5;
scale(1535) <= bm_5;
scale(1536) <= bm_5;
scale(1537) <= bm_5;
scale(1538) <= r;
scale(1539) <= f_4;
scale(1540) <= f_4;
scale(1541) <= f_4;
scale(1542) <= r;
scale(1543) <= g_4;
scale(1544) <= g_4;
scale(1545) <= g_4;
scale(1546) <= r;
scale(1547) <= a_5;
scale(1548) <= a_5;
scale(1549) <= a_5;
scale(1550) <= a_5;
----------------------end

led <= st;

piezo <= p_clk;
piezo2<= p_clk2;
--------------------------------------------------piezo1
process(clk,rst,rss)
begin
  if rst = '1' or rss = '1' then
	  cnt <= 0;
  elsif clk'event and clk = '1' and st = '1' then
     if cnt >= scale(note) then
	     cnt <= 0;
	  else
	     cnt <= cnt + 1;
	  end if;
  end if;
end process;


process (clk,rss,rst)
begin
if rss = '1' or rst = '1' then
  p_clk <= '0';
elsif clk'event and clk = '1' then
	if cnt = 1 then
		p_clk <= not p_clk;
	end if;
end if;
end process;
------------------------------------------------piezo2
process(clk,rst,rss)
begin
  if rst = '1' or rss = '1' then
	  cnt2 <= 0;
  elsif clk'event and clk = '1' and st = '1' then
     if cnt2 >= scale2(note) then
	     cnt2 <= 0;
	  else
	     cnt2 <= cnt2 + 1;
	  end if;
  end if;
end process;


process (clk,rss,rst)
begin
if rss = '1' or rst = '1' then
  p_clk2 <= '0';
elsif clk'event and clk = '1' then
	if cnt2 = 1 then
		p_clk2 <= not p_clk2;
	end if;
end if;
end process;


end a;